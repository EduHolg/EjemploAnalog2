magic
tech sky130A
magscale 1 2
timestamp 1715220266
<< pwell >>
rect 2270 -584 4432 -536
<< viali >>
rect 1476 700 1611 755
rect 2549 700 4381 770
rect 1465 -688 1600 -633
rect 2552 -698 4384 -628
<< metal1 >>
rect 780 961 5116 1161
rect 979 544 1133 961
rect 1443 755 1643 961
rect 1443 700 1476 755
rect 1611 700 1643 755
rect 1443 683 1643 700
rect 979 384 1133 390
rect 1203 648 1247 651
rect 1203 604 1580 648
rect 1203 321 1247 604
rect 2100 570 2168 961
rect 2513 770 4415 961
rect 2513 700 2549 770
rect 4381 700 4415 770
rect 2513 686 4415 700
rect 2264 596 4426 644
rect 1316 390 1322 544
rect 1476 390 1524 544
rect 1558 384 1939 546
rect 2094 502 2100 570
rect 2168 502 2174 570
rect 1203 277 1578 321
rect 798 28 998 107
rect 1203 28 1247 277
rect 798 -16 1247 28
rect 798 -93 998 -16
rect 1203 -231 1247 -16
rect 1777 87 1939 384
rect 2264 312 2312 596
rect 2468 508 2478 566
rect 2538 508 2548 566
rect 2662 506 2672 564
rect 2732 506 2742 564
rect 2856 506 2866 564
rect 2926 506 2936 564
rect 3046 506 3056 564
rect 3116 506 3126 564
rect 3236 506 3246 564
rect 3306 506 3316 564
rect 3428 506 3438 564
rect 3498 506 3508 564
rect 3622 508 3632 566
rect 3692 508 3702 566
rect 3812 506 3822 564
rect 3882 506 3892 564
rect 4006 508 4016 566
rect 4076 508 4086 566
rect 4196 508 4206 566
rect 4266 508 4276 566
rect 4390 506 4400 564
rect 4460 506 4470 564
rect 2564 364 2574 422
rect 2634 364 2644 422
rect 2756 366 2766 424
rect 2826 366 2836 424
rect 2948 364 2958 422
rect 3018 364 3028 422
rect 3140 364 3150 422
rect 3210 364 3220 422
rect 3332 364 3342 422
rect 3402 364 3412 422
rect 3522 366 3532 424
rect 3592 366 3602 424
rect 3716 364 3726 422
rect 3786 364 3796 422
rect 3908 364 3918 422
rect 3978 364 3988 422
rect 4098 364 4108 422
rect 4168 364 4178 422
rect 4292 364 4302 422
rect 4362 364 4372 422
rect 4660 362 4666 430
rect 4734 362 4740 430
rect 2264 264 4430 312
rect 2264 87 2312 264
rect 1777 -75 2312 87
rect 4666 42 4734 362
rect 4915 42 5115 107
rect 4666 26 5115 42
rect 1203 -275 1565 -231
rect 975 -330 1133 -324
rect 975 -869 1133 -488
rect 1203 -539 1247 -275
rect 1777 -327 1939 -75
rect 1302 -488 1308 -330
rect 1466 -488 1510 -330
rect 1549 -489 1939 -327
rect 2264 -222 2312 -75
rect 4660 -26 5115 26
rect 4660 -28 4734 -26
rect 2264 -270 4432 -222
rect 2094 -496 2100 -428
rect 2168 -496 2174 -428
rect 1203 -583 1558 -539
rect 1431 -633 1631 -620
rect 1431 -688 1465 -633
rect 1600 -688 1631 -633
rect 1431 -869 1631 -688
rect 2100 -869 2168 -496
rect 2264 -536 2312 -270
rect 4660 -294 4728 -28
rect 4915 -93 5115 -26
rect 2546 -358 2556 -300
rect 2616 -358 2626 -300
rect 2736 -358 2746 -300
rect 2806 -358 2816 -300
rect 2930 -358 2940 -300
rect 3000 -358 3010 -300
rect 3120 -356 3130 -298
rect 3190 -356 3200 -298
rect 3314 -356 3324 -298
rect 3384 -356 3394 -298
rect 3506 -356 3516 -298
rect 3576 -356 3586 -298
rect 3698 -358 3708 -300
rect 3768 -358 3778 -300
rect 3890 -358 3900 -300
rect 3960 -358 3970 -300
rect 4082 -358 4092 -300
rect 4152 -358 4162 -300
rect 4274 -360 4284 -302
rect 4344 -360 4354 -302
rect 4654 -362 4660 -294
rect 4728 -362 4734 -294
rect 2448 -492 2458 -434
rect 2518 -492 2528 -434
rect 2640 -492 2650 -434
rect 2710 -492 2720 -434
rect 2834 -492 2844 -434
rect 2904 -492 2914 -434
rect 3024 -494 3034 -436
rect 3094 -494 3104 -436
rect 3218 -492 3228 -434
rect 3288 -492 3298 -434
rect 3408 -492 3418 -434
rect 3478 -492 3488 -434
rect 3600 -492 3610 -434
rect 3670 -492 3680 -434
rect 3794 -492 3804 -434
rect 3864 -492 3874 -434
rect 3984 -492 3994 -434
rect 4054 -492 4064 -434
rect 4180 -490 4190 -432
rect 4250 -490 4260 -432
rect 4370 -492 4380 -434
rect 4440 -492 4450 -434
rect 2264 -584 4432 -536
rect 2499 -628 4426 -614
rect 2499 -698 2552 -628
rect 4384 -698 4426 -628
rect 2499 -869 4426 -698
rect 792 -1069 5110 -869
<< via1 >>
rect 979 390 1133 544
rect 1322 390 1476 544
rect 2100 502 2168 570
rect 2478 508 2538 566
rect 2672 506 2732 564
rect 2866 506 2926 564
rect 3056 506 3116 564
rect 3246 506 3306 564
rect 3438 506 3498 564
rect 3632 508 3692 566
rect 3822 506 3882 564
rect 4016 508 4076 566
rect 4206 508 4266 566
rect 4400 506 4460 564
rect 2574 364 2634 422
rect 2766 366 2826 424
rect 2958 364 3018 422
rect 3150 364 3210 422
rect 3342 364 3402 422
rect 3532 366 3592 424
rect 3726 364 3786 422
rect 3918 364 3978 422
rect 4108 364 4168 422
rect 4302 364 4362 422
rect 4666 362 4734 430
rect 975 -488 1133 -330
rect 1308 -488 1466 -330
rect 2100 -496 2168 -428
rect 2556 -358 2616 -300
rect 2746 -358 2806 -300
rect 2940 -358 3000 -300
rect 3130 -356 3190 -298
rect 3324 -356 3384 -298
rect 3516 -356 3576 -298
rect 3708 -358 3768 -300
rect 3900 -358 3960 -300
rect 4092 -358 4152 -300
rect 4284 -360 4344 -302
rect 4660 -362 4728 -294
rect 2458 -492 2518 -434
rect 2650 -492 2710 -434
rect 2844 -492 2904 -434
rect 3034 -494 3094 -436
rect 3228 -492 3288 -434
rect 3418 -492 3478 -434
rect 3610 -492 3670 -434
rect 3804 -492 3864 -434
rect 3994 -492 4054 -434
rect 4190 -490 4250 -432
rect 4380 -492 4440 -434
<< metal2 >>
rect 2100 570 2168 576
rect 2478 570 2538 576
rect 2672 570 2732 574
rect 2866 570 2926 574
rect 3056 570 3116 574
rect 3246 570 3306 574
rect 3438 570 3498 574
rect 3632 570 3692 576
rect 3822 570 3882 574
rect 4016 570 4076 576
rect 4206 570 4266 576
rect 4400 570 4460 574
rect 1322 544 1476 550
rect 973 390 979 544
rect 1133 390 1322 544
rect 2168 566 4492 570
rect 2168 508 2478 566
rect 2538 564 3632 566
rect 2538 508 2672 564
rect 2168 506 2672 508
rect 2732 506 2866 564
rect 2926 506 3056 564
rect 3116 506 3246 564
rect 3306 506 3438 564
rect 3498 508 3632 564
rect 3692 564 4016 566
rect 3692 508 3822 564
rect 3498 506 3822 508
rect 3882 508 4016 564
rect 4076 508 4206 566
rect 4266 564 4492 566
rect 4266 508 4400 564
rect 3882 506 4400 508
rect 4460 506 4492 564
rect 2168 502 4492 506
rect 2100 496 2168 502
rect 2478 498 2538 502
rect 2672 496 2732 502
rect 2866 496 2926 502
rect 3056 496 3116 502
rect 3246 496 3306 502
rect 3438 496 3498 502
rect 3632 498 3692 502
rect 3822 496 3882 502
rect 4016 498 4076 502
rect 4206 498 4266 502
rect 4400 496 4460 502
rect 2574 430 2634 432
rect 2766 430 2826 434
rect 2958 430 3018 432
rect 3150 430 3210 432
rect 3342 430 3402 432
rect 3532 430 3592 434
rect 3726 430 3786 432
rect 3918 430 3978 432
rect 4108 430 4168 432
rect 4302 430 4362 432
rect 4666 430 4734 436
rect 1322 384 1476 390
rect 2098 424 4666 430
rect 2098 422 2766 424
rect 2098 364 2574 422
rect 2634 366 2766 422
rect 2826 422 3532 424
rect 2826 366 2958 422
rect 2634 364 2958 366
rect 3018 364 3150 422
rect 3210 364 3342 422
rect 3402 366 3532 422
rect 3592 422 4666 424
rect 3592 366 3726 422
rect 3402 364 3726 366
rect 3786 364 3918 422
rect 3978 364 4108 422
rect 4168 364 4302 422
rect 4362 364 4666 422
rect 2098 362 4666 364
rect 2574 354 2634 362
rect 2766 356 2826 362
rect 2958 354 3018 362
rect 3150 354 3210 362
rect 3342 354 3402 362
rect 3532 356 3592 362
rect 3726 354 3786 362
rect 3918 354 3978 362
rect 4108 354 4168 362
rect 4302 354 4362 362
rect 4666 356 4734 362
rect 2556 -294 2616 -290
rect 2746 -294 2806 -290
rect 2940 -294 3000 -290
rect 3130 -294 3190 -288
rect 3324 -294 3384 -288
rect 3516 -294 3576 -288
rect 3708 -294 3768 -290
rect 3900 -294 3960 -290
rect 4092 -294 4152 -290
rect 4284 -294 4344 -292
rect 4660 -294 4728 -288
rect 2100 -298 4660 -294
rect 2100 -300 3130 -298
rect 1308 -330 1466 -324
rect 969 -488 975 -330
rect 1133 -488 1308 -330
rect 2100 -358 2556 -300
rect 2616 -358 2746 -300
rect 2806 -358 2940 -300
rect 3000 -356 3130 -300
rect 3190 -356 3324 -298
rect 3384 -356 3516 -298
rect 3576 -300 4660 -298
rect 3576 -356 3708 -300
rect 3000 -358 3708 -356
rect 3768 -358 3900 -300
rect 3960 -358 4092 -300
rect 4152 -302 4660 -300
rect 4152 -358 4284 -302
rect 2100 -360 4284 -358
rect 4344 -360 4660 -302
rect 2100 -362 4660 -360
rect 2556 -368 2616 -362
rect 2746 -368 2806 -362
rect 2940 -368 3000 -362
rect 3130 -366 3190 -362
rect 3324 -366 3384 -362
rect 3516 -366 3576 -362
rect 3708 -368 3768 -362
rect 3900 -368 3960 -362
rect 4092 -368 4152 -362
rect 4284 -370 4344 -362
rect 4660 -368 4728 -362
rect 1308 -494 1466 -488
rect 2100 -428 2168 -422
rect 2458 -428 2518 -424
rect 2650 -428 2710 -424
rect 2844 -428 2904 -424
rect 3034 -428 3094 -426
rect 3228 -428 3288 -424
rect 3418 -428 3478 -424
rect 3610 -428 3670 -424
rect 3804 -428 3864 -424
rect 3994 -428 4054 -424
rect 4190 -428 4250 -422
rect 4380 -428 4440 -424
rect 2168 -432 4492 -428
rect 2168 -434 4190 -432
rect 2168 -492 2458 -434
rect 2518 -492 2650 -434
rect 2710 -492 2844 -434
rect 2904 -436 3228 -434
rect 2904 -492 3034 -436
rect 2168 -494 3034 -492
rect 3094 -492 3228 -436
rect 3288 -492 3418 -434
rect 3478 -492 3610 -434
rect 3670 -492 3804 -434
rect 3864 -492 3994 -434
rect 4054 -490 4190 -434
rect 4250 -434 4492 -432
rect 4250 -490 4380 -434
rect 4054 -492 4380 -490
rect 4440 -492 4492 -434
rect 3094 -494 4492 -492
rect 2168 -496 4492 -494
rect 2100 -502 2168 -496
rect 2458 -502 2518 -496
rect 2650 -502 2710 -496
rect 2844 -502 2904 -496
rect 3034 -504 3094 -496
rect 3228 -502 3288 -496
rect 3418 -502 3478 -496
rect 3610 -502 3670 -496
rect 3804 -502 3864 -496
rect 3994 -502 4054 -496
rect 4190 -500 4250 -496
rect 4380 -502 4440 -496
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1715209795
transform 1 0 1543 0 1 463
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1715209795
transform 1 0 1529 0 1 -406
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_YTLFGX  XM3
timestamp 1715209795
transform 1 0 3449 0 1 -399
box -1127 -310 1127 310
use sky130_fd_pr__pfet_01v8_8DVCWJ  XM4
timestamp 1715209795
transform 1 0 3469 0 1 457
box -1127 -319 1127 319
<< labels >>
flabel metal1 780 961 980 1161 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 792 -1069 992 -869 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 798 -93 998 107 0 FreeSans 256 0 0 0 IN
port 3 nsew
flabel metal1 4915 -93 5115 107 0 FreeSans 256 0 0 0 OUT
port 2 nsew
<< end >>
