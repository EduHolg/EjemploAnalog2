magic
tech sky130A
magscale 1 2
timestamp 1717016881
<< nwell >>
rect -496 -279 496 279
<< pmos >>
rect -300 -60 300 60
<< pdiff >>
rect -358 17 -300 60
rect -358 -17 -346 17
rect -312 -17 -300 17
rect -358 -60 -300 -17
rect 300 17 358 60
rect 300 -17 312 17
rect 346 -17 358 17
rect 300 -60 358 -17
<< pdiffc >>
rect -346 -17 -312 17
rect 312 -17 346 17
<< nsubdiff >>
rect -460 209 -357 243
rect -323 209 -289 243
rect -255 209 -221 243
rect -187 209 -153 243
rect -119 209 -85 243
rect -51 209 -17 243
rect 17 209 51 243
rect 85 209 119 243
rect 153 209 187 243
rect 221 209 255 243
rect 289 209 323 243
rect 357 209 460 243
rect -460 119 -426 209
rect -460 51 -426 85
rect 426 119 460 209
rect -460 -17 -426 17
rect -460 -85 -426 -51
rect 426 51 460 85
rect 426 -17 460 17
rect -460 -209 -426 -119
rect 426 -85 460 -51
rect 426 -209 460 -119
rect -460 -243 -357 -209
rect -323 -243 -289 -209
rect -255 -243 -221 -209
rect -187 -243 -153 -209
rect -119 -243 -85 -209
rect -51 -243 -17 -209
rect 17 -243 51 -209
rect 85 -243 119 -209
rect 153 -243 187 -209
rect 221 -243 255 -209
rect 289 -243 323 -209
rect 357 -243 460 -209
<< nsubdiffcont >>
rect -357 209 -323 243
rect -289 209 -255 243
rect -221 209 -187 243
rect -153 209 -119 243
rect -85 209 -51 243
rect -17 209 17 243
rect 51 209 85 243
rect 119 209 153 243
rect 187 209 221 243
rect 255 209 289 243
rect 323 209 357 243
rect -460 85 -426 119
rect 426 85 460 119
rect -460 17 -426 51
rect -460 -51 -426 -17
rect 426 17 460 51
rect 426 -51 460 -17
rect -460 -119 -426 -85
rect 426 -119 460 -85
rect -357 -243 -323 -209
rect -289 -243 -255 -209
rect -221 -243 -187 -209
rect -153 -243 -119 -209
rect -85 -243 -51 -209
rect -17 -243 17 -209
rect 51 -243 85 -209
rect 119 -243 153 -209
rect 187 -243 221 -209
rect 255 -243 289 -209
rect 323 -243 357 -209
<< poly >>
rect -300 141 300 157
rect -300 107 -255 141
rect -221 107 -187 141
rect -153 107 -119 141
rect -85 107 -51 141
rect -17 107 17 141
rect 51 107 85 141
rect 119 107 153 141
rect 187 107 221 141
rect 255 107 300 141
rect -300 60 300 107
rect -300 -107 300 -60
rect -300 -141 -255 -107
rect -221 -141 -187 -107
rect -153 -141 -119 -107
rect -85 -141 -51 -107
rect -17 -141 17 -107
rect 51 -141 85 -107
rect 119 -141 153 -107
rect 187 -141 221 -107
rect 255 -141 300 -107
rect -300 -157 300 -141
<< polycont >>
rect -255 107 -221 141
rect -187 107 -153 141
rect -119 107 -85 141
rect -51 107 -17 141
rect 17 107 51 141
rect 85 107 119 141
rect 153 107 187 141
rect 221 107 255 141
rect -255 -141 -221 -107
rect -187 -141 -153 -107
rect -119 -141 -85 -107
rect -51 -141 -17 -107
rect 17 -141 51 -107
rect 85 -141 119 -107
rect 153 -141 187 -107
rect 221 -141 255 -107
<< locali >>
rect -460 209 -357 243
rect -323 209 -289 243
rect -255 209 -221 243
rect -187 209 -153 243
rect -119 209 -85 243
rect -51 209 -17 243
rect 17 209 51 243
rect 85 209 119 243
rect 153 209 187 243
rect 221 209 255 243
rect 289 209 323 243
rect 357 209 460 243
rect -460 119 -426 209
rect -300 107 -269 141
rect -221 107 -197 141
rect -153 107 -125 141
rect -85 107 -53 141
rect -17 107 17 141
rect 53 107 85 141
rect 125 107 153 141
rect 197 107 221 141
rect 269 107 300 141
rect 426 119 460 209
rect -460 51 -426 85
rect -460 -17 -426 17
rect -460 -85 -426 -51
rect -346 17 -312 64
rect -346 -64 -312 -17
rect 312 17 346 64
rect 312 -64 346 -17
rect 426 51 460 85
rect 426 -17 460 17
rect 426 -85 460 -51
rect -460 -209 -426 -119
rect -300 -141 -269 -107
rect -221 -141 -197 -107
rect -153 -141 -125 -107
rect -85 -141 -53 -107
rect -17 -141 17 -107
rect 53 -141 85 -107
rect 125 -141 153 -107
rect 197 -141 221 -107
rect 269 -141 300 -107
rect 426 -209 460 -119
rect -460 -243 -357 -209
rect -323 -243 -289 -209
rect -255 -243 -221 -209
rect -187 -243 -153 -209
rect -119 -243 -85 -209
rect -51 -243 -17 -209
rect 17 -243 51 -209
rect 85 -243 119 -209
rect 153 -243 187 -209
rect 221 -243 255 -209
rect 289 -243 323 -209
rect 357 -243 460 -209
<< viali >>
rect -269 107 -255 141
rect -255 107 -235 141
rect -197 107 -187 141
rect -187 107 -163 141
rect -125 107 -119 141
rect -119 107 -91 141
rect -53 107 -51 141
rect -51 107 -19 141
rect 19 107 51 141
rect 51 107 53 141
rect 91 107 119 141
rect 119 107 125 141
rect 163 107 187 141
rect 187 107 197 141
rect 235 107 255 141
rect 255 107 269 141
rect -346 -17 -312 17
rect 312 -17 346 17
rect -269 -141 -255 -107
rect -255 -141 -235 -107
rect -197 -141 -187 -107
rect -187 -141 -163 -107
rect -125 -141 -119 -107
rect -119 -141 -91 -107
rect -53 -141 -51 -107
rect -51 -141 -19 -107
rect 19 -141 51 -107
rect 51 -141 53 -107
rect 91 -141 119 -107
rect 119 -141 125 -107
rect 163 -141 187 -107
rect 187 -141 197 -107
rect 235 -141 255 -107
rect 255 -141 269 -107
<< metal1 >>
rect -296 141 296 147
rect -296 107 -269 141
rect -235 107 -197 141
rect -163 107 -125 141
rect -91 107 -53 141
rect -19 107 19 141
rect 53 107 91 141
rect 125 107 163 141
rect 197 107 235 141
rect 269 107 296 141
rect -296 101 296 107
rect -352 17 -306 60
rect -352 -17 -346 17
rect -312 -17 -306 17
rect -352 -60 -306 -17
rect 306 17 352 60
rect 306 -17 312 17
rect 346 -17 352 17
rect 306 -60 352 -17
rect -296 -107 296 -101
rect -296 -141 -269 -107
rect -235 -141 -197 -107
rect -163 -141 -125 -107
rect -91 -141 -53 -107
rect -19 -141 19 -107
rect 53 -141 91 -107
rect 125 -141 163 -107
rect 197 -141 235 -107
rect 269 -141 296 -107
rect -296 -147 296 -141
<< properties >>
string FIXED_BBOX -443 -226 443 226
<< end >>
