magic
tech sky130A
magscale 1 2
timestamp 1717016881
<< nwell >>
rect -496 -519 496 519
<< pmos >>
rect -300 -300 300 300
<< pdiff >>
rect -358 255 -300 300
rect -358 221 -346 255
rect -312 221 -300 255
rect -358 187 -300 221
rect -358 153 -346 187
rect -312 153 -300 187
rect -358 119 -300 153
rect -358 85 -346 119
rect -312 85 -300 119
rect -358 51 -300 85
rect -358 17 -346 51
rect -312 17 -300 51
rect -358 -17 -300 17
rect -358 -51 -346 -17
rect -312 -51 -300 -17
rect -358 -85 -300 -51
rect -358 -119 -346 -85
rect -312 -119 -300 -85
rect -358 -153 -300 -119
rect -358 -187 -346 -153
rect -312 -187 -300 -153
rect -358 -221 -300 -187
rect -358 -255 -346 -221
rect -312 -255 -300 -221
rect -358 -300 -300 -255
rect 300 255 358 300
rect 300 221 312 255
rect 346 221 358 255
rect 300 187 358 221
rect 300 153 312 187
rect 346 153 358 187
rect 300 119 358 153
rect 300 85 312 119
rect 346 85 358 119
rect 300 51 358 85
rect 300 17 312 51
rect 346 17 358 51
rect 300 -17 358 17
rect 300 -51 312 -17
rect 346 -51 358 -17
rect 300 -85 358 -51
rect 300 -119 312 -85
rect 346 -119 358 -85
rect 300 -153 358 -119
rect 300 -187 312 -153
rect 346 -187 358 -153
rect 300 -221 358 -187
rect 300 -255 312 -221
rect 346 -255 358 -221
rect 300 -300 358 -255
<< pdiffc >>
rect -346 221 -312 255
rect -346 153 -312 187
rect -346 85 -312 119
rect -346 17 -312 51
rect -346 -51 -312 -17
rect -346 -119 -312 -85
rect -346 -187 -312 -153
rect -346 -255 -312 -221
rect 312 221 346 255
rect 312 153 346 187
rect 312 85 346 119
rect 312 17 346 51
rect 312 -51 346 -17
rect 312 -119 346 -85
rect 312 -187 346 -153
rect 312 -255 346 -221
<< nsubdiff >>
rect -460 449 -357 483
rect -323 449 -289 483
rect -255 449 -221 483
rect -187 449 -153 483
rect -119 449 -85 483
rect -51 449 -17 483
rect 17 449 51 483
rect 85 449 119 483
rect 153 449 187 483
rect 221 449 255 483
rect 289 449 323 483
rect 357 449 460 483
rect -460 357 -426 449
rect -460 289 -426 323
rect 426 357 460 449
rect -460 221 -426 255
rect -460 153 -426 187
rect -460 85 -426 119
rect -460 17 -426 51
rect -460 -51 -426 -17
rect -460 -119 -426 -85
rect -460 -187 -426 -153
rect -460 -255 -426 -221
rect -460 -323 -426 -289
rect 426 289 460 323
rect 426 221 460 255
rect 426 153 460 187
rect 426 85 460 119
rect 426 17 460 51
rect 426 -51 460 -17
rect 426 -119 460 -85
rect 426 -187 460 -153
rect 426 -255 460 -221
rect -460 -449 -426 -357
rect 426 -323 460 -289
rect 426 -449 460 -357
rect -460 -483 -357 -449
rect -323 -483 -289 -449
rect -255 -483 -221 -449
rect -187 -483 -153 -449
rect -119 -483 -85 -449
rect -51 -483 -17 -449
rect 17 -483 51 -449
rect 85 -483 119 -449
rect 153 -483 187 -449
rect 221 -483 255 -449
rect 289 -483 323 -449
rect 357 -483 460 -449
<< nsubdiffcont >>
rect -357 449 -323 483
rect -289 449 -255 483
rect -221 449 -187 483
rect -153 449 -119 483
rect -85 449 -51 483
rect -17 449 17 483
rect 51 449 85 483
rect 119 449 153 483
rect 187 449 221 483
rect 255 449 289 483
rect 323 449 357 483
rect -460 323 -426 357
rect 426 323 460 357
rect -460 255 -426 289
rect -460 187 -426 221
rect -460 119 -426 153
rect -460 51 -426 85
rect -460 -17 -426 17
rect -460 -85 -426 -51
rect -460 -153 -426 -119
rect -460 -221 -426 -187
rect -460 -289 -426 -255
rect 426 255 460 289
rect 426 187 460 221
rect 426 119 460 153
rect 426 51 460 85
rect 426 -17 460 17
rect 426 -85 460 -51
rect 426 -153 460 -119
rect 426 -221 460 -187
rect 426 -289 460 -255
rect -460 -357 -426 -323
rect 426 -357 460 -323
rect -357 -483 -323 -449
rect -289 -483 -255 -449
rect -221 -483 -187 -449
rect -153 -483 -119 -449
rect -85 -483 -51 -449
rect -17 -483 17 -449
rect 51 -483 85 -449
rect 119 -483 153 -449
rect 187 -483 221 -449
rect 255 -483 289 -449
rect 323 -483 357 -449
<< poly >>
rect -300 381 300 397
rect -300 347 -255 381
rect -221 347 -187 381
rect -153 347 -119 381
rect -85 347 -51 381
rect -17 347 17 381
rect 51 347 85 381
rect 119 347 153 381
rect 187 347 221 381
rect 255 347 300 381
rect -300 300 300 347
rect -300 -347 300 -300
rect -300 -381 -255 -347
rect -221 -381 -187 -347
rect -153 -381 -119 -347
rect -85 -381 -51 -347
rect -17 -381 17 -347
rect 51 -381 85 -347
rect 119 -381 153 -347
rect 187 -381 221 -347
rect 255 -381 300 -347
rect -300 -397 300 -381
<< polycont >>
rect -255 347 -221 381
rect -187 347 -153 381
rect -119 347 -85 381
rect -51 347 -17 381
rect 17 347 51 381
rect 85 347 119 381
rect 153 347 187 381
rect 221 347 255 381
rect -255 -381 -221 -347
rect -187 -381 -153 -347
rect -119 -381 -85 -347
rect -51 -381 -17 -347
rect 17 -381 51 -347
rect 85 -381 119 -347
rect 153 -381 187 -347
rect 221 -381 255 -347
<< locali >>
rect -460 449 -357 483
rect -323 449 -289 483
rect -255 449 -221 483
rect -187 449 -153 483
rect -119 449 -85 483
rect -51 449 -17 483
rect 17 449 51 483
rect 85 449 119 483
rect 153 449 187 483
rect 221 449 255 483
rect 289 449 323 483
rect 357 449 460 483
rect -460 357 -426 449
rect -300 347 -269 381
rect -221 347 -197 381
rect -153 347 -125 381
rect -85 347 -53 381
rect -17 347 17 381
rect 53 347 85 381
rect 125 347 153 381
rect 197 347 221 381
rect 269 347 300 381
rect 426 357 460 449
rect -460 289 -426 323
rect -460 221 -426 255
rect -460 153 -426 187
rect -460 85 -426 119
rect -460 17 -426 51
rect -460 -51 -426 -17
rect -460 -119 -426 -85
rect -460 -187 -426 -153
rect -460 -255 -426 -221
rect -460 -323 -426 -289
rect -346 269 -312 304
rect -346 197 -312 221
rect -346 125 -312 153
rect -346 53 -312 85
rect -346 -17 -312 17
rect -346 -85 -312 -53
rect -346 -153 -312 -125
rect -346 -221 -312 -197
rect -346 -304 -312 -269
rect 312 269 346 304
rect 312 197 346 221
rect 312 125 346 153
rect 312 53 346 85
rect 312 -17 346 17
rect 312 -85 346 -53
rect 312 -153 346 -125
rect 312 -221 346 -197
rect 312 -304 346 -269
rect 426 289 460 323
rect 426 221 460 255
rect 426 153 460 187
rect 426 85 460 119
rect 426 17 460 51
rect 426 -51 460 -17
rect 426 -119 460 -85
rect 426 -187 460 -153
rect 426 -255 460 -221
rect 426 -323 460 -289
rect -460 -449 -426 -357
rect -300 -381 -269 -347
rect -221 -381 -197 -347
rect -153 -381 -125 -347
rect -85 -381 -53 -347
rect -17 -381 17 -347
rect 53 -381 85 -347
rect 125 -381 153 -347
rect 197 -381 221 -347
rect 269 -381 300 -347
rect 426 -449 460 -357
rect -460 -483 -357 -449
rect -323 -483 -289 -449
rect -255 -483 -221 -449
rect -187 -483 -153 -449
rect -119 -483 -85 -449
rect -51 -483 -17 -449
rect 17 -483 51 -449
rect 85 -483 119 -449
rect 153 -483 187 -449
rect 221 -483 255 -449
rect 289 -483 323 -449
rect 357 -483 460 -449
<< viali >>
rect -269 347 -255 381
rect -255 347 -235 381
rect -197 347 -187 381
rect -187 347 -163 381
rect -125 347 -119 381
rect -119 347 -91 381
rect -53 347 -51 381
rect -51 347 -19 381
rect 19 347 51 381
rect 51 347 53 381
rect 91 347 119 381
rect 119 347 125 381
rect 163 347 187 381
rect 187 347 197 381
rect 235 347 255 381
rect 255 347 269 381
rect -346 255 -312 269
rect -346 235 -312 255
rect -346 187 -312 197
rect -346 163 -312 187
rect -346 119 -312 125
rect -346 91 -312 119
rect -346 51 -312 53
rect -346 19 -312 51
rect -346 -51 -312 -19
rect -346 -53 -312 -51
rect -346 -119 -312 -91
rect -346 -125 -312 -119
rect -346 -187 -312 -163
rect -346 -197 -312 -187
rect -346 -255 -312 -235
rect -346 -269 -312 -255
rect 312 255 346 269
rect 312 235 346 255
rect 312 187 346 197
rect 312 163 346 187
rect 312 119 346 125
rect 312 91 346 119
rect 312 51 346 53
rect 312 19 346 51
rect 312 -51 346 -19
rect 312 -53 346 -51
rect 312 -119 346 -91
rect 312 -125 346 -119
rect 312 -187 346 -163
rect 312 -197 346 -187
rect 312 -255 346 -235
rect 312 -269 346 -255
rect -269 -381 -255 -347
rect -255 -381 -235 -347
rect -197 -381 -187 -347
rect -187 -381 -163 -347
rect -125 -381 -119 -347
rect -119 -381 -91 -347
rect -53 -381 -51 -347
rect -51 -381 -19 -347
rect 19 -381 51 -347
rect 51 -381 53 -347
rect 91 -381 119 -347
rect 119 -381 125 -347
rect 163 -381 187 -347
rect 187 -381 197 -347
rect 235 -381 255 -347
rect 255 -381 269 -347
<< metal1 >>
rect -296 381 296 387
rect -296 347 -269 381
rect -235 347 -197 381
rect -163 347 -125 381
rect -91 347 -53 381
rect -19 347 19 381
rect 53 347 91 381
rect 125 347 163 381
rect 197 347 235 381
rect 269 347 296 381
rect -296 341 296 347
rect -352 269 -306 300
rect -352 235 -346 269
rect -312 235 -306 269
rect -352 197 -306 235
rect -352 163 -346 197
rect -312 163 -306 197
rect -352 125 -306 163
rect -352 91 -346 125
rect -312 91 -306 125
rect -352 53 -306 91
rect -352 19 -346 53
rect -312 19 -306 53
rect -352 -19 -306 19
rect -352 -53 -346 -19
rect -312 -53 -306 -19
rect -352 -91 -306 -53
rect -352 -125 -346 -91
rect -312 -125 -306 -91
rect -352 -163 -306 -125
rect -352 -197 -346 -163
rect -312 -197 -306 -163
rect -352 -235 -306 -197
rect -352 -269 -346 -235
rect -312 -269 -306 -235
rect -352 -300 -306 -269
rect 306 269 352 300
rect 306 235 312 269
rect 346 235 352 269
rect 306 197 352 235
rect 306 163 312 197
rect 346 163 352 197
rect 306 125 352 163
rect 306 91 312 125
rect 346 91 352 125
rect 306 53 352 91
rect 306 19 312 53
rect 346 19 352 53
rect 306 -19 352 19
rect 306 -53 312 -19
rect 346 -53 352 -19
rect 306 -91 352 -53
rect 306 -125 312 -91
rect 346 -125 352 -91
rect 306 -163 352 -125
rect 306 -197 312 -163
rect 346 -197 352 -163
rect 306 -235 352 -197
rect 306 -269 312 -235
rect 346 -269 352 -235
rect 306 -300 352 -269
rect -296 -347 296 -341
rect -296 -381 -269 -347
rect -235 -381 -197 -347
rect -163 -381 -125 -347
rect -91 -381 -53 -347
rect -19 -381 19 -347
rect 53 -381 91 -347
rect 125 -381 163 -347
rect 197 -381 235 -347
rect 269 -381 296 -347
rect -296 -387 296 -381
<< properties >>
string FIXED_BBOX -443 -466 443 466
<< end >>
