magic
tech sky130A
magscale 1 2
timestamp 1717016881
<< pwell >>
rect -686 -500 686 500
<< nmos >>
rect -500 -300 500 300
<< ndiff >>
rect -558 255 -500 300
rect -558 221 -546 255
rect -512 221 -500 255
rect -558 187 -500 221
rect -558 153 -546 187
rect -512 153 -500 187
rect -558 119 -500 153
rect -558 85 -546 119
rect -512 85 -500 119
rect -558 51 -500 85
rect -558 17 -546 51
rect -512 17 -500 51
rect -558 -17 -500 17
rect -558 -51 -546 -17
rect -512 -51 -500 -17
rect -558 -85 -500 -51
rect -558 -119 -546 -85
rect -512 -119 -500 -85
rect -558 -153 -500 -119
rect -558 -187 -546 -153
rect -512 -187 -500 -153
rect -558 -221 -500 -187
rect -558 -255 -546 -221
rect -512 -255 -500 -221
rect -558 -300 -500 -255
rect 500 255 558 300
rect 500 221 512 255
rect 546 221 558 255
rect 500 187 558 221
rect 500 153 512 187
rect 546 153 558 187
rect 500 119 558 153
rect 500 85 512 119
rect 546 85 558 119
rect 500 51 558 85
rect 500 17 512 51
rect 546 17 558 51
rect 500 -17 558 17
rect 500 -51 512 -17
rect 546 -51 558 -17
rect 500 -85 558 -51
rect 500 -119 512 -85
rect 546 -119 558 -85
rect 500 -153 558 -119
rect 500 -187 512 -153
rect 546 -187 558 -153
rect 500 -221 558 -187
rect 500 -255 512 -221
rect 546 -255 558 -221
rect 500 -300 558 -255
<< ndiffc >>
rect -546 221 -512 255
rect -546 153 -512 187
rect -546 85 -512 119
rect -546 17 -512 51
rect -546 -51 -512 -17
rect -546 -119 -512 -85
rect -546 -187 -512 -153
rect -546 -255 -512 -221
rect 512 221 546 255
rect 512 153 546 187
rect 512 85 546 119
rect 512 17 546 51
rect 512 -51 546 -17
rect 512 -119 546 -85
rect 512 -187 546 -153
rect 512 -255 546 -221
<< psubdiff >>
rect -660 440 -561 474
rect -527 440 -493 474
rect -459 440 -425 474
rect -391 440 -357 474
rect -323 440 -289 474
rect -255 440 -221 474
rect -187 440 -153 474
rect -119 440 -85 474
rect -51 440 -17 474
rect 17 440 51 474
rect 85 440 119 474
rect 153 440 187 474
rect 221 440 255 474
rect 289 440 323 474
rect 357 440 391 474
rect 425 440 459 474
rect 493 440 527 474
rect 561 440 660 474
rect -660 357 -626 440
rect -660 289 -626 323
rect 626 357 660 440
rect -660 221 -626 255
rect -660 153 -626 187
rect -660 85 -626 119
rect -660 17 -626 51
rect -660 -51 -626 -17
rect -660 -119 -626 -85
rect -660 -187 -626 -153
rect -660 -255 -626 -221
rect -660 -323 -626 -289
rect 626 289 660 323
rect 626 221 660 255
rect 626 153 660 187
rect 626 85 660 119
rect 626 17 660 51
rect 626 -51 660 -17
rect 626 -119 660 -85
rect 626 -187 660 -153
rect 626 -255 660 -221
rect -660 -440 -626 -357
rect 626 -323 660 -289
rect 626 -440 660 -357
rect -660 -474 -561 -440
rect -527 -474 -493 -440
rect -459 -474 -425 -440
rect -391 -474 -357 -440
rect -323 -474 -289 -440
rect -255 -474 -221 -440
rect -187 -474 -153 -440
rect -119 -474 -85 -440
rect -51 -474 -17 -440
rect 17 -474 51 -440
rect 85 -474 119 -440
rect 153 -474 187 -440
rect 221 -474 255 -440
rect 289 -474 323 -440
rect 357 -474 391 -440
rect 425 -474 459 -440
rect 493 -474 527 -440
rect 561 -474 660 -440
<< psubdiffcont >>
rect -561 440 -527 474
rect -493 440 -459 474
rect -425 440 -391 474
rect -357 440 -323 474
rect -289 440 -255 474
rect -221 440 -187 474
rect -153 440 -119 474
rect -85 440 -51 474
rect -17 440 17 474
rect 51 440 85 474
rect 119 440 153 474
rect 187 440 221 474
rect 255 440 289 474
rect 323 440 357 474
rect 391 440 425 474
rect 459 440 493 474
rect 527 440 561 474
rect -660 323 -626 357
rect 626 323 660 357
rect -660 255 -626 289
rect -660 187 -626 221
rect -660 119 -626 153
rect -660 51 -626 85
rect -660 -17 -626 17
rect -660 -85 -626 -51
rect -660 -153 -626 -119
rect -660 -221 -626 -187
rect -660 -289 -626 -255
rect 626 255 660 289
rect 626 187 660 221
rect 626 119 660 153
rect 626 51 660 85
rect 626 -17 660 17
rect 626 -85 660 -51
rect 626 -153 660 -119
rect 626 -221 660 -187
rect 626 -289 660 -255
rect -660 -357 -626 -323
rect 626 -357 660 -323
rect -561 -474 -527 -440
rect -493 -474 -459 -440
rect -425 -474 -391 -440
rect -357 -474 -323 -440
rect -289 -474 -255 -440
rect -221 -474 -187 -440
rect -153 -474 -119 -440
rect -85 -474 -51 -440
rect -17 -474 17 -440
rect 51 -474 85 -440
rect 119 -474 153 -440
rect 187 -474 221 -440
rect 255 -474 289 -440
rect 323 -474 357 -440
rect 391 -474 425 -440
rect 459 -474 493 -440
rect 527 -474 561 -440
<< poly >>
rect -500 372 500 388
rect -500 338 -459 372
rect -425 338 -391 372
rect -357 338 -323 372
rect -289 338 -255 372
rect -221 338 -187 372
rect -153 338 -119 372
rect -85 338 -51 372
rect -17 338 17 372
rect 51 338 85 372
rect 119 338 153 372
rect 187 338 221 372
rect 255 338 289 372
rect 323 338 357 372
rect 391 338 425 372
rect 459 338 500 372
rect -500 300 500 338
rect -500 -338 500 -300
rect -500 -372 -459 -338
rect -425 -372 -391 -338
rect -357 -372 -323 -338
rect -289 -372 -255 -338
rect -221 -372 -187 -338
rect -153 -372 -119 -338
rect -85 -372 -51 -338
rect -17 -372 17 -338
rect 51 -372 85 -338
rect 119 -372 153 -338
rect 187 -372 221 -338
rect 255 -372 289 -338
rect 323 -372 357 -338
rect 391 -372 425 -338
rect 459 -372 500 -338
rect -500 -388 500 -372
<< polycont >>
rect -459 338 -425 372
rect -391 338 -357 372
rect -323 338 -289 372
rect -255 338 -221 372
rect -187 338 -153 372
rect -119 338 -85 372
rect -51 338 -17 372
rect 17 338 51 372
rect 85 338 119 372
rect 153 338 187 372
rect 221 338 255 372
rect 289 338 323 372
rect 357 338 391 372
rect 425 338 459 372
rect -459 -372 -425 -338
rect -391 -372 -357 -338
rect -323 -372 -289 -338
rect -255 -372 -221 -338
rect -187 -372 -153 -338
rect -119 -372 -85 -338
rect -51 -372 -17 -338
rect 17 -372 51 -338
rect 85 -372 119 -338
rect 153 -372 187 -338
rect 221 -372 255 -338
rect 289 -372 323 -338
rect 357 -372 391 -338
rect 425 -372 459 -338
<< locali >>
rect -660 440 -561 474
rect -527 440 -493 474
rect -459 440 -425 474
rect -391 440 -357 474
rect -323 440 -289 474
rect -255 440 -221 474
rect -187 440 -153 474
rect -119 440 -85 474
rect -51 440 -17 474
rect 17 440 51 474
rect 85 440 119 474
rect 153 440 187 474
rect 221 440 255 474
rect 289 440 323 474
rect 357 440 391 474
rect 425 440 459 474
rect 493 440 527 474
rect 561 440 660 474
rect -660 357 -626 440
rect -500 338 -459 372
rect -415 338 -391 372
rect -343 338 -323 372
rect -271 338 -255 372
rect -199 338 -187 372
rect -127 338 -119 372
rect -55 338 -51 372
rect 51 338 55 372
rect 119 338 127 372
rect 187 338 199 372
rect 255 338 271 372
rect 323 338 343 372
rect 391 338 415 372
rect 459 338 500 372
rect 626 357 660 440
rect -660 289 -626 323
rect -660 221 -626 255
rect -660 153 -626 187
rect -660 85 -626 119
rect -660 17 -626 51
rect -660 -51 -626 -17
rect -660 -119 -626 -85
rect -660 -187 -626 -153
rect -660 -255 -626 -221
rect -660 -323 -626 -289
rect -546 269 -512 304
rect -546 197 -512 221
rect -546 125 -512 153
rect -546 53 -512 85
rect -546 -17 -512 17
rect -546 -85 -512 -53
rect -546 -153 -512 -125
rect -546 -221 -512 -197
rect -546 -304 -512 -269
rect 512 269 546 304
rect 512 197 546 221
rect 512 125 546 153
rect 512 53 546 85
rect 512 -17 546 17
rect 512 -85 546 -53
rect 512 -153 546 -125
rect 512 -221 546 -197
rect 512 -304 546 -269
rect 626 289 660 323
rect 626 221 660 255
rect 626 153 660 187
rect 626 85 660 119
rect 626 17 660 51
rect 626 -51 660 -17
rect 626 -119 660 -85
rect 626 -187 660 -153
rect 626 -255 660 -221
rect 626 -323 660 -289
rect -660 -440 -626 -357
rect -500 -372 -459 -338
rect -415 -372 -391 -338
rect -343 -372 -323 -338
rect -271 -372 -255 -338
rect -199 -372 -187 -338
rect -127 -372 -119 -338
rect -55 -372 -51 -338
rect 51 -372 55 -338
rect 119 -372 127 -338
rect 187 -372 199 -338
rect 255 -372 271 -338
rect 323 -372 343 -338
rect 391 -372 415 -338
rect 459 -372 500 -338
rect 626 -440 660 -357
rect -660 -474 -561 -440
rect -527 -474 -493 -440
rect -459 -474 -425 -440
rect -391 -474 -357 -440
rect -323 -474 -289 -440
rect -255 -474 -221 -440
rect -187 -474 -153 -440
rect -119 -474 -85 -440
rect -51 -474 -17 -440
rect 17 -474 51 -440
rect 85 -474 119 -440
rect 153 -474 187 -440
rect 221 -474 255 -440
rect 289 -474 323 -440
rect 357 -474 391 -440
rect 425 -474 459 -440
rect 493 -474 527 -440
rect 561 -474 660 -440
<< viali >>
rect -449 338 -425 372
rect -425 338 -415 372
rect -377 338 -357 372
rect -357 338 -343 372
rect -305 338 -289 372
rect -289 338 -271 372
rect -233 338 -221 372
rect -221 338 -199 372
rect -161 338 -153 372
rect -153 338 -127 372
rect -89 338 -85 372
rect -85 338 -55 372
rect -17 338 17 372
rect 55 338 85 372
rect 85 338 89 372
rect 127 338 153 372
rect 153 338 161 372
rect 199 338 221 372
rect 221 338 233 372
rect 271 338 289 372
rect 289 338 305 372
rect 343 338 357 372
rect 357 338 377 372
rect 415 338 425 372
rect 425 338 449 372
rect -546 255 -512 269
rect -546 235 -512 255
rect -546 187 -512 197
rect -546 163 -512 187
rect -546 119 -512 125
rect -546 91 -512 119
rect -546 51 -512 53
rect -546 19 -512 51
rect -546 -51 -512 -19
rect -546 -53 -512 -51
rect -546 -119 -512 -91
rect -546 -125 -512 -119
rect -546 -187 -512 -163
rect -546 -197 -512 -187
rect -546 -255 -512 -235
rect -546 -269 -512 -255
rect 512 255 546 269
rect 512 235 546 255
rect 512 187 546 197
rect 512 163 546 187
rect 512 119 546 125
rect 512 91 546 119
rect 512 51 546 53
rect 512 19 546 51
rect 512 -51 546 -19
rect 512 -53 546 -51
rect 512 -119 546 -91
rect 512 -125 546 -119
rect 512 -187 546 -163
rect 512 -197 546 -187
rect 512 -255 546 -235
rect 512 -269 546 -255
rect -449 -372 -425 -338
rect -425 -372 -415 -338
rect -377 -372 -357 -338
rect -357 -372 -343 -338
rect -305 -372 -289 -338
rect -289 -372 -271 -338
rect -233 -372 -221 -338
rect -221 -372 -199 -338
rect -161 -372 -153 -338
rect -153 -372 -127 -338
rect -89 -372 -85 -338
rect -85 -372 -55 -338
rect -17 -372 17 -338
rect 55 -372 85 -338
rect 85 -372 89 -338
rect 127 -372 153 -338
rect 153 -372 161 -338
rect 199 -372 221 -338
rect 221 -372 233 -338
rect 271 -372 289 -338
rect 289 -372 305 -338
rect 343 -372 357 -338
rect 357 -372 377 -338
rect 415 -372 425 -338
rect 425 -372 449 -338
<< metal1 >>
rect -496 372 496 378
rect -496 338 -449 372
rect -415 338 -377 372
rect -343 338 -305 372
rect -271 338 -233 372
rect -199 338 -161 372
rect -127 338 -89 372
rect -55 338 -17 372
rect 17 338 55 372
rect 89 338 127 372
rect 161 338 199 372
rect 233 338 271 372
rect 305 338 343 372
rect 377 338 415 372
rect 449 338 496 372
rect -496 332 496 338
rect -552 269 -506 300
rect -552 235 -546 269
rect -512 235 -506 269
rect -552 197 -506 235
rect -552 163 -546 197
rect -512 163 -506 197
rect -552 125 -506 163
rect -552 91 -546 125
rect -512 91 -506 125
rect -552 53 -506 91
rect -552 19 -546 53
rect -512 19 -506 53
rect -552 -19 -506 19
rect -552 -53 -546 -19
rect -512 -53 -506 -19
rect -552 -91 -506 -53
rect -552 -125 -546 -91
rect -512 -125 -506 -91
rect -552 -163 -506 -125
rect -552 -197 -546 -163
rect -512 -197 -506 -163
rect -552 -235 -506 -197
rect -552 -269 -546 -235
rect -512 -269 -506 -235
rect -552 -300 -506 -269
rect 506 269 552 300
rect 506 235 512 269
rect 546 235 552 269
rect 506 197 552 235
rect 506 163 512 197
rect 546 163 552 197
rect 506 125 552 163
rect 506 91 512 125
rect 546 91 552 125
rect 506 53 552 91
rect 506 19 512 53
rect 546 19 552 53
rect 506 -19 552 19
rect 506 -53 512 -19
rect 546 -53 552 -19
rect 506 -91 552 -53
rect 506 -125 512 -91
rect 546 -125 552 -91
rect 506 -163 552 -125
rect 506 -197 512 -163
rect 546 -197 552 -163
rect 506 -235 552 -197
rect 506 -269 512 -235
rect 546 -269 552 -235
rect 506 -300 552 -269
rect -496 -338 496 -332
rect -496 -372 -449 -338
rect -415 -372 -377 -338
rect -343 -372 -305 -338
rect -271 -372 -233 -338
rect -199 -372 -161 -338
rect -127 -372 -89 -338
rect -55 -372 -17 -338
rect 17 -372 55 -338
rect 89 -372 127 -338
rect 161 -372 199 -338
rect 233 -372 271 -338
rect 305 -372 343 -338
rect 377 -372 415 -338
rect 449 -372 496 -338
rect -496 -378 496 -372
<< properties >>
string FIXED_BBOX -642 -456 642 456
<< end >>
