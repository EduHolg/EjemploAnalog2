magic
tech sky130A
magscale 1 2
timestamp 1717016881
<< locali >>
rect 8036 1022 8080 1032
rect 8036 988 8041 1022
rect 8075 988 8080 1022
rect 13684 1010 13730 1032
rect 8036 950 8080 988
rect 8036 916 8041 950
rect 8075 916 8080 950
rect 8036 878 8080 916
rect 8036 844 8041 878
rect 8075 844 8080 878
rect 8036 806 8080 844
rect 8036 772 8041 806
rect 8075 772 8080 806
rect 7220 763 7610 768
rect 7220 729 7254 763
rect 7288 729 7326 763
rect 7360 729 7398 763
rect 7432 729 7470 763
rect 7504 729 7542 763
rect 7576 729 7610 763
rect 7220 724 7610 729
rect 8036 734 8080 772
rect 11134 994 11178 1004
rect 11134 960 11139 994
rect 11173 960 11178 994
rect 11134 922 11178 960
rect 11134 888 11139 922
rect 11173 888 11178 922
rect 11134 850 11178 888
rect 11134 816 11139 850
rect 11173 816 11178 850
rect 11134 778 11178 816
rect 11134 744 11139 778
rect 11173 744 11178 778
rect 11134 734 11178 744
rect 12420 994 12468 1004
rect 12420 960 12427 994
rect 12461 960 12468 994
rect 12420 922 12468 960
rect 12420 888 12427 922
rect 12461 888 12468 922
rect 12420 850 12468 888
rect 12420 816 12427 850
rect 12461 816 12468 850
rect 12420 778 12468 816
rect 12420 744 12427 778
rect 12461 744 12468 778
rect 12420 734 12468 744
rect 13684 976 13690 1010
rect 13724 976 13730 1010
rect 13684 938 13730 976
rect 13684 904 13690 938
rect 13724 904 13730 938
rect 13684 866 13730 904
rect 13684 832 13690 866
rect 13724 832 13730 866
rect 13684 794 13730 832
rect 13684 760 13690 794
rect 13724 760 13730 794
rect 13684 738 13730 760
rect 14208 764 14596 768
rect 8036 700 8041 734
rect 8075 700 8080 734
rect 14208 730 14241 764
rect 14275 730 14313 764
rect 14347 730 14385 764
rect 14419 730 14457 764
rect 14491 730 14529 764
rect 14563 730 14596 764
rect 14208 726 14596 730
rect 8036 662 8080 700
rect 8036 628 8041 662
rect 8075 628 8080 662
rect 8036 590 8080 628
rect 8036 556 8041 590
rect 8075 556 8080 590
rect 8036 518 8080 556
rect 8036 484 8041 518
rect 8075 484 8080 518
rect 8036 446 8080 484
rect 8036 412 8041 446
rect 8075 412 8080 446
rect 8036 374 8080 412
rect 8036 340 8041 374
rect 8075 340 8080 374
rect 8036 302 8080 340
rect 8036 268 8041 302
rect 8075 268 8080 302
rect 8036 258 8080 268
rect 12794 206 12840 216
rect 12794 172 12800 206
rect 12834 172 12840 206
rect 12794 134 12840 172
rect 12794 100 12800 134
rect 12834 100 12840 134
rect 12794 62 12840 100
rect 12794 28 12800 62
rect 12834 28 12840 62
rect 12794 -10 12840 28
rect 12794 -44 12800 -10
rect 12834 -44 12840 -10
rect 12794 -82 12840 -44
rect 12794 -116 12800 -82
rect 12834 -116 12840 -82
rect 12794 -154 12840 -116
rect 12794 -188 12800 -154
rect 12834 -188 12840 -154
rect 12794 -226 12840 -188
rect 12794 -260 12800 -226
rect 12834 -260 12840 -226
rect 8038 -271 8082 -260
rect 8038 -305 8043 -271
rect 8077 -305 8082 -271
rect 8038 -343 8082 -305
rect 8038 -377 8043 -343
rect 8077 -377 8082 -343
rect 8038 -415 8082 -377
rect 8038 -449 8043 -415
rect 8077 -449 8082 -415
rect 8038 -487 8082 -449
rect 8038 -521 8043 -487
rect 8077 -521 8082 -487
rect 8038 -559 8082 -521
rect 8038 -593 8043 -559
rect 8077 -593 8082 -559
rect 8038 -631 8082 -593
rect 8038 -665 8043 -631
rect 8077 -665 8082 -631
rect 8038 -703 8082 -665
rect 8038 -737 8043 -703
rect 8077 -737 8082 -703
rect 8038 -775 8082 -737
rect 8038 -809 8043 -775
rect 8077 -809 8082 -775
rect 8038 -847 8082 -809
rect 8038 -881 8043 -847
rect 8077 -881 8082 -847
rect 8038 -919 8082 -881
rect 8038 -953 8043 -919
rect 8077 -953 8082 -919
rect 8038 -991 8082 -953
rect 8038 -1025 8043 -991
rect 8077 -1025 8082 -991
rect 8038 -1036 8082 -1025
rect 8926 -271 8968 -260
rect 8926 -305 8930 -271
rect 8964 -305 8968 -271
rect 8926 -343 8968 -305
rect 8926 -377 8930 -343
rect 8964 -377 8968 -343
rect 8926 -415 8968 -377
rect 8926 -449 8930 -415
rect 8964 -449 8968 -415
rect 8926 -487 8968 -449
rect 8926 -521 8930 -487
rect 8964 -521 8968 -487
rect 8926 -559 8968 -521
rect 12794 -298 12840 -260
rect 12794 -332 12800 -298
rect 12834 -332 12840 -298
rect 12794 -370 12840 -332
rect 12794 -404 12800 -370
rect 12834 -404 12840 -370
rect 12794 -442 12840 -404
rect 12794 -476 12800 -442
rect 12834 -476 12840 -442
rect 12794 -514 12840 -476
rect 12794 -548 12800 -514
rect 12834 -548 12840 -514
rect 12794 -558 12840 -548
rect 13680 206 13726 216
rect 13680 172 13686 206
rect 13720 172 13726 206
rect 13680 134 13726 172
rect 13680 100 13686 134
rect 13720 100 13726 134
rect 13680 62 13726 100
rect 13680 28 13686 62
rect 13720 28 13726 62
rect 13680 -10 13726 28
rect 13680 -44 13686 -10
rect 13720 -44 13726 -10
rect 13680 -82 13726 -44
rect 13680 -116 13686 -82
rect 13720 -116 13726 -82
rect 13680 -154 13726 -116
rect 13680 -188 13686 -154
rect 13720 -188 13726 -154
rect 13680 -226 13726 -188
rect 13680 -260 13686 -226
rect 13720 -260 13726 -226
rect 13680 -298 13726 -260
rect 13680 -332 13686 -298
rect 13720 -332 13726 -298
rect 13680 -370 13726 -332
rect 13680 -404 13686 -370
rect 13720 -404 13726 -370
rect 13680 -442 13726 -404
rect 13680 -476 13686 -442
rect 13720 -476 13726 -442
rect 13680 -514 13726 -476
rect 13680 -548 13686 -514
rect 13720 -548 13726 -514
rect 13680 -558 13726 -548
rect 8926 -593 8930 -559
rect 8964 -593 8968 -559
rect 8926 -631 8968 -593
rect 8926 -665 8930 -631
rect 8964 -665 8968 -631
rect 8926 -703 8968 -665
rect 8926 -737 8930 -703
rect 8964 -737 8968 -703
rect 8926 -775 8968 -737
rect 8926 -809 8930 -775
rect 8964 -809 8968 -775
rect 8926 -847 8968 -809
rect 8926 -881 8930 -847
rect 8964 -881 8968 -847
rect 8926 -919 8968 -881
rect 8926 -953 8930 -919
rect 8964 -953 8968 -919
rect 8926 -991 8968 -953
rect 8926 -1025 8930 -991
rect 8964 -1025 8968 -991
rect 8926 -1036 8968 -1025
rect 12796 -1088 12842 -1078
rect 11132 -1099 11176 -1098
rect 11132 -1133 11137 -1099
rect 11171 -1133 11176 -1099
rect 11132 -1171 11176 -1133
rect 11132 -1205 11137 -1171
rect 11171 -1205 11176 -1171
rect 11132 -1243 11176 -1205
rect 11132 -1277 11137 -1243
rect 11171 -1277 11176 -1243
rect 11132 -1315 11176 -1277
rect 11132 -1349 11137 -1315
rect 11171 -1349 11176 -1315
rect 11132 -1387 11176 -1349
rect 11132 -1421 11137 -1387
rect 11171 -1421 11176 -1387
rect 11132 -1459 11176 -1421
rect 11132 -1493 11137 -1459
rect 11171 -1493 11176 -1459
rect 11132 -1531 11176 -1493
rect 8036 -1578 8080 -1556
rect 8036 -1612 8041 -1578
rect 8075 -1612 8080 -1578
rect 8036 -1650 8080 -1612
rect 8036 -1684 8041 -1650
rect 8075 -1684 8080 -1650
rect 8036 -1722 8080 -1684
rect 8036 -1756 8041 -1722
rect 8075 -1756 8080 -1722
rect 8036 -1794 8080 -1756
rect 8036 -1828 8041 -1794
rect 8075 -1828 8080 -1794
rect 8036 -1850 8080 -1828
rect 8922 -1578 8966 -1556
rect 8922 -1612 8927 -1578
rect 8961 -1612 8966 -1578
rect 11132 -1565 11137 -1531
rect 11171 -1565 11176 -1531
rect 8922 -1650 8966 -1612
rect 8922 -1684 8927 -1650
rect 8961 -1684 8966 -1650
rect 8922 -1722 8966 -1684
rect 8922 -1756 8927 -1722
rect 8961 -1756 8966 -1722
rect 8922 -1794 8966 -1756
rect 8922 -1828 8927 -1794
rect 8961 -1828 8966 -1794
rect 8922 -1850 8966 -1828
rect 9322 -1592 9374 -1582
rect 9322 -1626 9331 -1592
rect 9365 -1626 9374 -1592
rect 9322 -1664 9374 -1626
rect 9322 -1698 9331 -1664
rect 9365 -1698 9374 -1664
rect 9322 -1736 9374 -1698
rect 9322 -1770 9331 -1736
rect 9365 -1770 9374 -1736
rect 9322 -1808 9374 -1770
rect 9322 -1842 9331 -1808
rect 9365 -1842 9374 -1808
rect 9322 -1852 9374 -1842
rect 10612 -1592 10660 -1582
rect 10612 -1626 10619 -1592
rect 10653 -1626 10660 -1592
rect 10612 -1664 10660 -1626
rect 10612 -1698 10619 -1664
rect 10653 -1698 10660 -1664
rect 10612 -1736 10660 -1698
rect 10612 -1770 10619 -1736
rect 10653 -1770 10660 -1736
rect 10612 -1808 10660 -1770
rect 10612 -1842 10619 -1808
rect 10653 -1842 10660 -1808
rect 10612 -1852 10660 -1842
rect 11132 -1603 11176 -1565
rect 11132 -1637 11137 -1603
rect 11171 -1637 11176 -1603
rect 11132 -1675 11176 -1637
rect 11132 -1709 11137 -1675
rect 11171 -1709 11176 -1675
rect 11132 -1747 11176 -1709
rect 11132 -1781 11137 -1747
rect 11171 -1781 11176 -1747
rect 11132 -1819 11176 -1781
rect 11132 -1853 11137 -1819
rect 11171 -1853 11176 -1819
rect 12796 -1122 12802 -1088
rect 12836 -1122 12842 -1088
rect 12796 -1160 12842 -1122
rect 12796 -1194 12802 -1160
rect 12836 -1194 12842 -1160
rect 12796 -1232 12842 -1194
rect 12796 -1266 12802 -1232
rect 12836 -1266 12842 -1232
rect 12796 -1304 12842 -1266
rect 12796 -1338 12802 -1304
rect 12836 -1338 12842 -1304
rect 12796 -1376 12842 -1338
rect 12796 -1410 12802 -1376
rect 12836 -1410 12842 -1376
rect 12796 -1448 12842 -1410
rect 12796 -1482 12802 -1448
rect 12836 -1482 12842 -1448
rect 12796 -1520 12842 -1482
rect 12796 -1554 12802 -1520
rect 12836 -1554 12842 -1520
rect 12796 -1592 12842 -1554
rect 12796 -1626 12802 -1592
rect 12836 -1626 12842 -1592
rect 12796 -1664 12842 -1626
rect 12796 -1698 12802 -1664
rect 12836 -1698 12842 -1664
rect 12796 -1736 12842 -1698
rect 12796 -1770 12802 -1736
rect 12836 -1770 12842 -1736
rect 12796 -1808 12842 -1770
rect 12796 -1842 12802 -1808
rect 12836 -1842 12842 -1808
rect 12796 -1852 12842 -1842
rect 13684 -1088 13726 -1078
rect 13684 -1122 13688 -1088
rect 13722 -1122 13726 -1088
rect 13684 -1160 13726 -1122
rect 13684 -1194 13688 -1160
rect 13722 -1194 13726 -1160
rect 13684 -1232 13726 -1194
rect 13684 -1266 13688 -1232
rect 13722 -1266 13726 -1232
rect 13684 -1304 13726 -1266
rect 13684 -1338 13688 -1304
rect 13722 -1338 13726 -1304
rect 13684 -1376 13726 -1338
rect 13684 -1410 13688 -1376
rect 13722 -1410 13726 -1376
rect 13684 -1448 13726 -1410
rect 13684 -1482 13688 -1448
rect 13722 -1482 13726 -1448
rect 13684 -1520 13726 -1482
rect 13684 -1554 13688 -1520
rect 13722 -1554 13726 -1520
rect 13684 -1592 13726 -1554
rect 13684 -1626 13688 -1592
rect 13722 -1626 13726 -1592
rect 13684 -1664 13726 -1626
rect 13684 -1698 13688 -1664
rect 13722 -1698 13726 -1664
rect 13684 -1736 13726 -1698
rect 13684 -1770 13688 -1736
rect 13722 -1770 13726 -1736
rect 13684 -1808 13726 -1770
rect 13684 -1842 13688 -1808
rect 13722 -1842 13726 -1808
rect 13684 -1852 13726 -1842
rect 11132 -1854 11176 -1853
<< viali >>
rect 8041 988 8075 1022
rect 8041 916 8075 950
rect 8041 844 8075 878
rect 8041 772 8075 806
rect 7254 729 7288 763
rect 7326 729 7360 763
rect 7398 729 7432 763
rect 7470 729 7504 763
rect 7542 729 7576 763
rect 11139 960 11173 994
rect 11139 888 11173 922
rect 11139 816 11173 850
rect 11139 744 11173 778
rect 12427 960 12461 994
rect 12427 888 12461 922
rect 12427 816 12461 850
rect 12427 744 12461 778
rect 13690 976 13724 1010
rect 13690 904 13724 938
rect 13690 832 13724 866
rect 13690 760 13724 794
rect 8041 700 8075 734
rect 14241 730 14275 764
rect 14313 730 14347 764
rect 14385 730 14419 764
rect 14457 730 14491 764
rect 14529 730 14563 764
rect 8041 628 8075 662
rect 8041 556 8075 590
rect 8041 484 8075 518
rect 8041 412 8075 446
rect 8041 340 8075 374
rect 8041 268 8075 302
rect 12800 172 12834 206
rect 12800 100 12834 134
rect 12800 28 12834 62
rect 12800 -44 12834 -10
rect 12800 -116 12834 -82
rect 12800 -188 12834 -154
rect 12800 -260 12834 -226
rect 8043 -305 8077 -271
rect 8043 -377 8077 -343
rect 8043 -449 8077 -415
rect 8043 -521 8077 -487
rect 8043 -593 8077 -559
rect 8043 -665 8077 -631
rect 8043 -737 8077 -703
rect 8043 -809 8077 -775
rect 8043 -881 8077 -847
rect 8043 -953 8077 -919
rect 8043 -1025 8077 -991
rect 8930 -305 8964 -271
rect 8930 -377 8964 -343
rect 8930 -449 8964 -415
rect 8930 -521 8964 -487
rect 12800 -332 12834 -298
rect 12800 -404 12834 -370
rect 12800 -476 12834 -442
rect 12800 -548 12834 -514
rect 13686 172 13720 206
rect 13686 100 13720 134
rect 13686 28 13720 62
rect 13686 -44 13720 -10
rect 13686 -116 13720 -82
rect 13686 -188 13720 -154
rect 13686 -260 13720 -226
rect 13686 -332 13720 -298
rect 13686 -404 13720 -370
rect 13686 -476 13720 -442
rect 13686 -548 13720 -514
rect 8930 -593 8964 -559
rect 8930 -665 8964 -631
rect 8930 -737 8964 -703
rect 8930 -809 8964 -775
rect 8930 -881 8964 -847
rect 8930 -953 8964 -919
rect 8930 -1025 8964 -991
rect 11137 -1133 11171 -1099
rect 11137 -1205 11171 -1171
rect 11137 -1277 11171 -1243
rect 11137 -1349 11171 -1315
rect 11137 -1421 11171 -1387
rect 11137 -1493 11171 -1459
rect 8041 -1612 8075 -1578
rect 8041 -1684 8075 -1650
rect 8041 -1756 8075 -1722
rect 8041 -1828 8075 -1794
rect 8927 -1612 8961 -1578
rect 11137 -1565 11171 -1531
rect 8927 -1684 8961 -1650
rect 8927 -1756 8961 -1722
rect 8927 -1828 8961 -1794
rect 9331 -1626 9365 -1592
rect 9331 -1698 9365 -1664
rect 9331 -1770 9365 -1736
rect 9331 -1842 9365 -1808
rect 10619 -1626 10653 -1592
rect 10619 -1698 10653 -1664
rect 10619 -1770 10653 -1736
rect 10619 -1842 10653 -1808
rect 11137 -1637 11171 -1603
rect 11137 -1709 11171 -1675
rect 11137 -1781 11171 -1747
rect 11137 -1853 11171 -1819
rect 12802 -1122 12836 -1088
rect 12802 -1194 12836 -1160
rect 12802 -1266 12836 -1232
rect 12802 -1338 12836 -1304
rect 12802 -1410 12836 -1376
rect 12802 -1482 12836 -1448
rect 12802 -1554 12836 -1520
rect 12802 -1626 12836 -1592
rect 12802 -1698 12836 -1664
rect 12802 -1770 12836 -1736
rect 12802 -1842 12836 -1808
rect 13688 -1122 13722 -1088
rect 13688 -1194 13722 -1160
rect 13688 -1266 13722 -1232
rect 13688 -1338 13722 -1304
rect 13688 -1410 13722 -1376
rect 13688 -1482 13722 -1448
rect 13688 -1554 13722 -1520
rect 13688 -1626 13722 -1592
rect 13688 -1698 13722 -1664
rect 13688 -1770 13722 -1736
rect 13688 -1842 13722 -1808
<< metal1 >>
rect 7096 1396 14726 1502
rect 8036 1140 8084 1396
rect 12326 1232 12938 1270
rect 8024 1022 8094 1140
rect 8024 988 8041 1022
rect 8075 988 8094 1022
rect 8024 950 8094 988
rect 8024 916 8041 950
rect 8075 916 8094 950
rect 8024 878 8094 916
rect 11122 994 11192 1116
rect 11122 960 11139 994
rect 11173 960 11192 994
rect 11122 922 11192 960
rect 11122 888 11139 922
rect 11173 888 11192 922
rect 12326 908 12370 1232
rect 12408 994 12484 1118
rect 12408 960 12427 994
rect 12461 960 12484 994
rect 12408 922 12484 960
rect 12408 888 12427 922
rect 12461 888 12484 922
rect 12894 908 12938 1232
rect 13690 1144 13738 1396
rect 13672 1010 13746 1144
rect 13672 976 13690 1010
rect 13724 976 13746 1010
rect 13672 938 13746 976
rect 13672 904 13690 938
rect 13724 904 13746 938
rect 13672 898 13746 904
rect 8024 844 8041 878
rect 8075 844 8094 878
rect 8024 806 8094 844
rect 10748 850 11266 888
rect 10748 826 11139 850
rect 7104 763 7726 788
rect 7104 729 7254 763
rect 7288 729 7326 763
rect 7360 729 7398 763
rect 7432 729 7470 763
rect 7504 729 7542 763
rect 7576 729 7726 763
rect 7104 712 7726 729
rect 8024 772 8041 806
rect 8075 772 8094 806
rect 8024 734 8094 772
rect 8024 700 8041 734
rect 8075 700 8094 734
rect 8024 670 8094 700
rect 11122 816 11139 826
rect 11173 826 11266 850
rect 12408 850 12484 888
rect 11173 816 11192 826
rect 11122 778 11192 816
rect 12408 816 12427 850
rect 12461 816 12484 850
rect 12958 836 12960 888
rect 13584 866 13746 898
rect 13584 856 13690 866
rect 11122 744 11139 778
rect 11173 744 11192 778
rect 7236 576 7296 664
rect 8024 662 8186 670
rect 8024 628 8041 662
rect 8075 628 8186 662
rect 8830 630 9376 682
rect 8024 624 8186 628
rect 11122 624 11192 744
rect 8024 590 8094 624
rect 8024 556 8041 590
rect 8075 556 8094 590
rect 8024 518 8094 556
rect 8024 484 8041 518
rect 8075 484 8094 518
rect 8024 446 8094 484
rect 8024 412 8041 446
rect 8075 412 8094 446
rect 8024 374 8094 412
rect 8024 340 8041 374
rect 8075 340 8094 374
rect 8024 302 8094 340
rect 8024 268 8041 302
rect 8075 268 8094 302
rect 8024 -271 8094 268
rect 8024 -305 8043 -271
rect 8077 -305 8094 -271
rect 8460 -282 8520 294
rect 10452 34 10520 150
rect 11340 34 11412 786
rect 12408 778 12484 816
rect 12408 744 12427 778
rect 12461 744 12484 778
rect 13672 832 13690 856
rect 13724 832 13746 866
rect 13672 794 13746 832
rect 12408 622 12484 744
rect 10452 -40 11412 34
rect 10452 -42 10520 -40
rect 8024 -343 8094 -305
rect 8024 -377 8043 -343
rect 8077 -377 8094 -343
rect 8024 -415 8094 -377
rect 8786 -396 8852 -264
rect 8914 -271 8978 -142
rect 8914 -305 8930 -271
rect 8964 -305 8978 -271
rect 8914 -343 8978 -305
rect 8914 -377 8930 -343
rect 8964 -377 8978 -343
rect 8024 -449 8043 -415
rect 8077 -449 8094 -415
rect 8024 -487 8094 -449
rect 8024 -521 8043 -487
rect 8077 -521 8094 -487
rect 8024 -559 8094 -521
rect 8024 -593 8043 -559
rect 8077 -593 8094 -559
rect 8024 -630 8094 -593
rect 8914 -415 8978 -377
rect 12418 -380 12472 622
rect 8914 -449 8930 -415
rect 8964 -449 8978 -415
rect 8914 -487 8978 -449
rect 8914 -521 8930 -487
rect 8964 -521 8978 -487
rect 8914 -559 8978 -521
rect 8914 -593 8930 -559
rect 8964 -593 8978 -559
rect 8024 -631 8182 -630
rect 8024 -665 8043 -631
rect 8077 -665 8182 -631
rect 8024 -674 8182 -665
rect 8914 -631 8978 -593
rect 8914 -665 8930 -631
rect 8964 -665 8978 -631
rect 8024 -703 8094 -674
rect 8024 -737 8043 -703
rect 8077 -737 8094 -703
rect 8024 -775 8094 -737
rect 8024 -809 8043 -775
rect 8077 -809 8094 -775
rect 8024 -847 8094 -809
rect 8024 -881 8043 -847
rect 8077 -881 8094 -847
rect 8024 -919 8094 -881
rect 8024 -953 8043 -919
rect 8077 -953 8094 -919
rect 8024 -991 8094 -953
rect 8024 -1025 8043 -991
rect 8077 -1025 8094 -991
rect 8914 -703 8978 -665
rect 8914 -737 8930 -703
rect 8964 -737 8978 -703
rect 8914 -775 8978 -737
rect 8914 -809 8930 -775
rect 8964 -809 8978 -775
rect 8914 -847 8978 -809
rect 8914 -881 8930 -847
rect 8964 -881 8978 -847
rect 8914 -919 8978 -881
rect 8914 -953 8930 -919
rect 8964 -953 8978 -919
rect 8914 -991 8978 -953
rect 8024 -1142 8094 -1025
rect 8460 -1294 8520 -1012
rect 7574 -1346 8520 -1294
rect 7218 -2198 7258 -1388
rect 8024 -1578 8094 -1450
rect 8024 -1612 8041 -1578
rect 8075 -1612 8094 -1578
rect 8460 -1588 8520 -1346
rect 8914 -1025 8930 -991
rect 8964 -1025 8978 -991
rect 8914 -1578 8978 -1025
rect 9316 -448 12472 -380
rect 12784 206 12856 332
rect 12784 172 12800 206
rect 12834 172 12856 206
rect 13202 198 13262 774
rect 13672 760 13690 794
rect 13724 760 13746 794
rect 13672 206 13746 760
rect 14100 764 14710 782
rect 14100 730 14241 764
rect 14275 730 14313 764
rect 14347 730 14385 764
rect 14419 730 14457 764
rect 14491 730 14529 764
rect 14563 730 14710 764
rect 14100 714 14710 730
rect 14522 570 14582 658
rect 12784 134 12856 172
rect 12784 100 12800 134
rect 12834 100 12856 134
rect 12784 62 12856 100
rect 12784 28 12800 62
rect 12834 28 12856 62
rect 12784 -10 12856 28
rect 12784 -44 12800 -10
rect 12834 -44 12856 -10
rect 12784 -82 12856 -44
rect 12784 -116 12800 -82
rect 12834 -116 12856 -82
rect 12784 -154 12856 -116
rect 12784 -188 12800 -154
rect 12834 -188 12856 -154
rect 13672 172 13686 206
rect 13720 172 13746 206
rect 13672 134 13746 172
rect 13672 100 13686 134
rect 13720 100 13746 134
rect 13672 62 13746 100
rect 13672 28 13686 62
rect 13720 28 13746 62
rect 13672 -10 13746 28
rect 13672 -44 13686 -10
rect 13720 -44 13746 -10
rect 13672 -82 13746 -44
rect 13672 -116 13686 -82
rect 13720 -116 13746 -82
rect 13672 -154 13746 -116
rect 13672 -156 13686 -154
rect 12784 -226 12856 -188
rect 13580 -188 13686 -156
rect 13720 -188 13746 -154
rect 13580 -196 13746 -188
rect 12784 -260 12800 -226
rect 12834 -260 12856 -226
rect 12784 -298 12856 -260
rect 12784 -332 12800 -298
rect 12834 -332 12856 -298
rect 12784 -370 12856 -332
rect 12784 -404 12800 -370
rect 12834 -404 12856 -370
rect 12784 -442 12856 -404
rect 13672 -226 13746 -196
rect 13672 -260 13686 -226
rect 13720 -260 13746 -226
rect 13672 -298 13746 -260
rect 13672 -332 13686 -298
rect 13720 -332 13746 -298
rect 13672 -370 13746 -332
rect 13672 -404 13686 -370
rect 13720 -404 13746 -370
rect 9316 -1470 9380 -448
rect 12784 -476 12800 -442
rect 12834 -476 12856 -442
rect 12784 -514 12856 -476
rect 12784 -548 12800 -514
rect 12834 -548 12856 -514
rect 12916 -548 12982 -416
rect 13672 -442 13746 -404
rect 13672 -476 13686 -442
rect 13720 -476 13746 -442
rect 13672 -514 13746 -476
rect 10440 -856 11400 -782
rect 8024 -1650 8094 -1612
rect 8024 -1684 8041 -1650
rect 8075 -1682 8094 -1650
rect 8914 -1612 8927 -1578
rect 8961 -1612 8978 -1578
rect 8914 -1650 8978 -1612
rect 8075 -1684 8176 -1682
rect 8024 -1722 8176 -1684
rect 8914 -1684 8927 -1650
rect 8961 -1684 8978 -1650
rect 8024 -1756 8041 -1722
rect 8075 -1724 8176 -1722
rect 8075 -1756 8094 -1724
rect 8024 -1794 8094 -1756
rect 8024 -1828 8041 -1794
rect 8075 -1828 8094 -1794
rect 8024 -1954 8094 -1828
rect 8826 -2016 8874 -1702
rect 8914 -1722 8978 -1684
rect 8914 -1756 8927 -1722
rect 8961 -1756 8978 -1722
rect 8914 -1794 8978 -1756
rect 8914 -1828 8927 -1794
rect 8961 -1828 8978 -1794
rect 8914 -1964 8978 -1828
rect 9306 -1592 9384 -1470
rect 9306 -1626 9331 -1592
rect 9365 -1626 9384 -1592
rect 10440 -1608 10512 -856
rect 11120 -1099 11184 -980
rect 11120 -1133 11137 -1099
rect 11171 -1133 11184 -1099
rect 11332 -1126 11400 -856
rect 12784 -1088 12856 -548
rect 11120 -1171 11184 -1133
rect 11120 -1205 11137 -1171
rect 11171 -1205 11184 -1171
rect 12272 -1198 12340 -1100
rect 12784 -1122 12802 -1088
rect 12836 -1122 12856 -1088
rect 13272 -812 13332 -526
rect 13672 -548 13686 -514
rect 13720 -548 13746 -514
rect 13672 -672 13746 -548
rect 13272 -864 14250 -812
rect 13272 -1102 13332 -864
rect 13674 -1088 13742 -966
rect 12784 -1160 12856 -1122
rect 12784 -1194 12802 -1160
rect 12836 -1194 12856 -1160
rect 11120 -1243 11184 -1205
rect 11120 -1277 11137 -1243
rect 11171 -1277 11184 -1243
rect 11120 -1315 11184 -1277
rect 11120 -1349 11137 -1315
rect 11171 -1349 11184 -1315
rect 11120 -1387 11184 -1349
rect 11120 -1421 11137 -1387
rect 11171 -1421 11184 -1387
rect 11120 -1459 11184 -1421
rect 10604 -1592 10678 -1470
rect 9306 -1664 9384 -1626
rect 9306 -1698 9331 -1664
rect 9365 -1698 9384 -1664
rect 10604 -1626 10619 -1592
rect 10653 -1626 10678 -1592
rect 10604 -1664 10678 -1626
rect 10604 -1680 10619 -1664
rect 9306 -1736 9384 -1698
rect 10522 -1698 10619 -1680
rect 10653 -1680 10678 -1664
rect 11120 -1493 11137 -1459
rect 11171 -1493 11184 -1459
rect 11120 -1531 11184 -1493
rect 11120 -1565 11137 -1531
rect 11171 -1565 11184 -1531
rect 11120 -1603 11184 -1565
rect 11120 -1637 11137 -1603
rect 11171 -1637 11184 -1603
rect 11120 -1675 11184 -1637
rect 11120 -1680 11137 -1675
rect 10653 -1698 11137 -1680
rect 9306 -1770 9331 -1736
rect 9365 -1770 9384 -1736
rect 9306 -1808 9384 -1770
rect 9306 -1842 9331 -1808
rect 9365 -1842 9384 -1808
rect 9306 -1962 9384 -1842
rect 9416 -2016 9464 -1702
rect 10522 -1709 11137 -1698
rect 11171 -1680 11184 -1675
rect 12784 -1232 12856 -1194
rect 12784 -1266 12802 -1232
rect 12836 -1266 12856 -1232
rect 12784 -1304 12856 -1266
rect 12784 -1338 12802 -1304
rect 12836 -1338 12856 -1304
rect 12784 -1376 12856 -1338
rect 12784 -1410 12802 -1376
rect 12836 -1410 12856 -1376
rect 12784 -1448 12856 -1410
rect 13674 -1122 13688 -1088
rect 13722 -1122 13742 -1088
rect 13674 -1160 13742 -1122
rect 13674 -1194 13688 -1160
rect 13722 -1194 13742 -1160
rect 13674 -1232 13742 -1194
rect 13674 -1266 13688 -1232
rect 13722 -1266 13742 -1232
rect 13674 -1304 13742 -1266
rect 13674 -1338 13688 -1304
rect 13722 -1338 13742 -1304
rect 13674 -1376 13742 -1338
rect 13674 -1410 13688 -1376
rect 13722 -1410 13742 -1376
rect 13674 -1446 13742 -1410
rect 12784 -1482 12802 -1448
rect 12836 -1482 12856 -1448
rect 12784 -1520 12856 -1482
rect 13582 -1448 13742 -1446
rect 13582 -1482 13688 -1448
rect 13722 -1482 13742 -1448
rect 13582 -1486 13742 -1482
rect 12784 -1554 12802 -1520
rect 12836 -1554 12856 -1520
rect 12784 -1592 12856 -1554
rect 12784 -1626 12802 -1592
rect 12836 -1626 12856 -1592
rect 12784 -1664 12856 -1626
rect 11171 -1709 11270 -1680
rect 10522 -1736 11270 -1709
rect 12784 -1698 12802 -1664
rect 12836 -1698 12856 -1664
rect 10522 -1742 10619 -1736
rect 10604 -1770 10619 -1742
rect 10653 -1742 11270 -1736
rect 10653 -1770 10678 -1742
rect 10604 -1808 10678 -1770
rect 10604 -1842 10619 -1808
rect 10653 -1842 10678 -1808
rect 10604 -1964 10678 -1842
rect 8826 -2068 9464 -2016
rect 10824 -2198 10916 -1742
rect 11120 -1747 11184 -1742
rect 11120 -1781 11137 -1747
rect 11171 -1781 11184 -1747
rect 11120 -1819 11184 -1781
rect 11120 -1853 11137 -1819
rect 11171 -1853 11184 -1819
rect 11120 -1962 11184 -1853
rect 12340 -2020 12384 -1726
rect 12784 -1736 12856 -1698
rect 13674 -1520 13742 -1486
rect 13674 -1554 13688 -1520
rect 13722 -1554 13742 -1520
rect 13674 -1592 13742 -1554
rect 13674 -1626 13688 -1592
rect 13722 -1626 13742 -1592
rect 13674 -1664 13742 -1626
rect 13674 -1698 13688 -1664
rect 13722 -1698 13742 -1664
rect 12784 -1770 12802 -1736
rect 12836 -1770 12856 -1736
rect 12784 -1808 12856 -1770
rect 12784 -1842 12802 -1808
rect 12836 -1842 12856 -1808
rect 12784 -1964 12856 -1842
rect 12892 -2020 12936 -1726
rect 13674 -1736 13742 -1698
rect 13674 -1770 13688 -1736
rect 13722 -1770 13742 -1736
rect 13674 -1808 13742 -1770
rect 13674 -1842 13688 -1808
rect 13722 -1842 13742 -1808
rect 13674 -1966 13742 -1842
rect 12340 -2072 12936 -2020
rect 14562 -2198 14602 -1386
rect 7096 -2304 14726 -2198
use sky130_fd_pr__nfet_01v8_HXU4AK  sky130_fd_pr__nfet_01v8_HXU4AK_0
timestamp 1717016881
transform 1 0 11800 0 1 869
box -686 -257 686 257
use sky130_fd_pr__nfet_01v8_HXU4AK  sky130_fd_pr__nfet_01v8_HXU4AK_1
timestamp 1717016881
transform 1 0 9992 0 1 -1717
box -686 -257 686 257
use sky130_fd_pr__nfet_01v8_MXF53G  sky130_fd_pr__nfet_01v8_MXF53G_0
timestamp 1717016881
transform 1 0 11796 0 1 -1476
box -686 -500 686 500
use sky130_fd_pr__nfet_01v8_MXF53G  sky130_fd_pr__nfet_01v8_MXF53G_1
timestamp 1717016881
transform 1 0 10062 0 1 650
box -686 -500 686 500
use sky130_fd_pr__pfet_01v8_GE7BQD  sky130_fd_pr__pfet_01v8_GE7BQD_0
timestamp 1717016881
transform 1 0 14402 0 1 -419
box -326 -1219 326 1219
use sky130_fd_pr__pfet_01v8_GE7BQD  sky130_fd_pr__pfet_01v8_GE7BQD_1
timestamp 1717016881
transform 1 0 7414 0 1 -419
box -326 -1219 326 1219
use sky130_fd_pr__pfet_01v8_KDYT8F  sky130_fd_pr__pfet_01v8_KDYT8F_0
timestamp 1717016881
transform 1 0 13264 0 1 885
box -496 -279 496 279
use sky130_fd_pr__pfet_01v8_KDYT8F  sky130_fd_pr__pfet_01v8_KDYT8F_1
timestamp 1717016881
transform 1 0 8500 0 1 -1703
box -496 -279 496 279
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_0
timestamp 1717016881
transform -1 0 13260 0 -1 -171
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_1
timestamp 1717016881
transform -1 0 13262 0 -1 -1465
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_2
timestamp 1717016881
transform -1 0 8502 0 -1 645
box -496 -519 496 519
use sky130_fd_pr__pfet_01v8_NXK9QA  sky130_fd_pr__pfet_01v8_NXK9QA_3
timestamp 1717016881
transform -1 0 8503 0 -1 -648
box -496 -519 496 519
<< end >>
