VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_adennen_inverter
  CLASS BLOCK ;
  FOREIGN tt_um_adennen_inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.892600 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.892600 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.339300 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 16.568199 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 111.890 16.830 115.150 29.020 ;
        RECT 116.480 25.650 121.440 30.840 ;
      LAYER pwell ;
        RECT 123.330 25.770 130.190 30.770 ;
        RECT 132.020 28.080 138.880 30.650 ;
      LAYER nwell ;
        RECT 140.290 28.050 145.250 30.840 ;
        RECT 116.485 19.185 121.445 24.375 ;
        RECT 140.270 21.570 145.230 26.760 ;
        RECT 116.470 15.110 121.430 17.900 ;
      LAYER pwell ;
        RECT 122.980 15.150 129.840 17.720 ;
        RECT 132.000 15.140 138.860 20.140 ;
      LAYER nwell ;
        RECT 140.280 15.100 145.240 20.290 ;
        RECT 146.830 16.830 150.090 29.020 ;
      LAYER li1 ;
        RECT 116.660 30.490 121.260 30.660 ;
        RECT 116.660 30.180 116.830 30.490 ;
        RECT 112.550 28.840 114.500 28.860 ;
        RECT 112.070 28.670 114.970 28.840 ;
        RECT 112.070 17.180 112.240 28.670 ;
        RECT 112.550 28.640 114.500 28.670 ;
        RECT 112.870 28.160 114.170 28.330 ;
        RECT 112.640 17.905 112.810 27.945 ;
        RECT 114.230 17.905 114.400 27.945 ;
        RECT 112.870 17.520 114.170 17.690 ;
        RECT 114.800 17.180 114.970 28.670 ;
        RECT 116.630 26.310 116.850 30.180 ;
        RECT 117.460 29.980 120.460 30.150 ;
        RECT 117.230 26.725 117.400 29.765 ;
        RECT 120.520 26.725 120.690 29.765 ;
        RECT 117.460 26.340 120.460 26.510 ;
        RECT 116.660 26.000 116.830 26.310 ;
        RECT 121.090 26.000 121.260 30.490 ;
        RECT 116.660 25.830 121.260 26.000 ;
        RECT 123.460 30.470 130.060 30.640 ;
        RECT 123.460 26.070 123.630 30.470 ;
        RECT 124.260 29.960 129.260 30.130 ;
        RECT 124.030 26.750 124.200 29.790 ;
        RECT 129.320 26.750 129.490 29.790 ;
        RECT 124.260 26.410 129.260 26.580 ;
        RECT 129.890 26.070 130.060 30.470 ;
        RECT 132.150 30.350 138.750 30.520 ;
        RECT 132.150 30.040 132.320 30.350 ;
        RECT 138.580 30.040 138.750 30.350 ;
        RECT 140.470 30.490 145.070 30.660 ;
        RECT 132.120 28.690 132.340 30.040 ;
        RECT 132.950 29.840 137.950 30.010 ;
        RECT 132.720 29.060 132.890 29.670 ;
        RECT 138.010 29.060 138.180 29.670 ;
        RECT 132.950 28.720 137.950 28.890 ;
        RECT 138.550 28.690 138.790 30.040 ;
        RECT 132.150 28.380 132.320 28.690 ;
        RECT 138.580 28.380 138.750 28.690 ;
        RECT 132.150 28.210 138.750 28.380 ;
        RECT 140.470 28.400 140.640 30.490 ;
        RECT 144.900 30.180 145.070 30.490 ;
        RECT 141.270 29.980 144.270 30.150 ;
        RECT 141.040 29.125 141.210 29.765 ;
        RECT 144.330 29.125 144.500 29.765 ;
        RECT 141.270 28.740 144.270 28.910 ;
        RECT 144.870 28.710 145.100 30.180 ;
        RECT 147.490 28.840 149.430 28.860 ;
        RECT 144.900 28.400 145.070 28.710 ;
        RECT 140.470 28.230 145.070 28.400 ;
        RECT 147.010 28.670 149.910 28.840 ;
        RECT 140.450 26.410 145.050 26.580 ;
        RECT 140.450 26.100 140.620 26.410 ;
        RECT 144.880 26.100 145.050 26.410 ;
        RECT 123.460 25.900 130.060 26.070 ;
        RECT 116.665 24.025 121.265 24.195 ;
        RECT 116.665 23.720 116.835 24.025 ;
        RECT 121.095 23.720 121.265 24.025 ;
        RECT 116.640 19.840 116.860 23.720 ;
        RECT 117.465 23.515 120.465 23.685 ;
        RECT 117.235 20.260 117.405 23.300 ;
        RECT 120.525 20.260 120.695 23.300 ;
        RECT 117.465 19.875 120.465 20.045 ;
        RECT 121.080 19.840 121.290 23.720 ;
        RECT 140.420 22.230 140.650 26.100 ;
        RECT 141.250 25.900 144.250 26.070 ;
        RECT 141.020 22.645 141.190 25.685 ;
        RECT 144.310 22.645 144.480 25.685 ;
        RECT 141.250 22.260 144.250 22.430 ;
        RECT 144.850 22.230 145.080 26.100 ;
        RECT 140.450 21.920 140.620 22.230 ;
        RECT 144.880 21.920 145.050 22.230 ;
        RECT 140.450 21.750 145.050 21.920 ;
        RECT 132.130 19.840 138.730 20.010 ;
        RECT 116.665 19.535 116.835 19.840 ;
        RECT 121.095 19.535 121.265 19.840 ;
        RECT 116.665 19.365 121.265 19.535 ;
        RECT 132.130 19.530 132.300 19.840 ;
        RECT 116.650 17.550 121.250 17.720 ;
        RECT 116.650 17.240 116.820 17.550 ;
        RECT 121.080 17.240 121.250 17.550 ;
        RECT 123.110 17.420 129.710 17.590 ;
        RECT 112.070 17.010 114.970 17.180 ;
        RECT 116.630 15.770 116.850 17.240 ;
        RECT 117.450 17.040 120.450 17.210 ;
        RECT 117.220 16.185 117.390 16.825 ;
        RECT 120.510 16.185 120.680 16.825 ;
        RECT 117.450 15.800 120.450 15.970 ;
        RECT 121.060 15.770 121.280 17.240 ;
        RECT 123.110 17.110 123.280 17.420 ;
        RECT 129.540 17.110 129.710 17.420 ;
        RECT 116.650 15.460 116.820 15.770 ;
        RECT 121.080 15.460 121.250 15.770 ;
        RECT 123.060 15.760 123.320 17.110 ;
        RECT 123.910 16.910 128.910 17.080 ;
        RECT 123.680 16.130 123.850 16.740 ;
        RECT 128.970 16.130 129.140 16.740 ;
        RECT 123.910 15.790 128.910 15.960 ;
        RECT 129.510 15.760 129.750 17.110 ;
        RECT 116.650 15.290 121.250 15.460 ;
        RECT 123.110 15.450 123.280 15.760 ;
        RECT 129.540 15.450 129.710 15.760 ;
        RECT 132.110 15.750 132.330 19.530 ;
        RECT 132.930 19.330 137.930 19.500 ;
        RECT 132.700 16.120 132.870 19.160 ;
        RECT 137.990 16.120 138.160 19.160 ;
        RECT 132.930 15.780 137.930 15.950 ;
        RECT 123.110 15.280 129.710 15.450 ;
        RECT 132.130 15.440 132.300 15.750 ;
        RECT 138.560 15.440 138.730 19.840 ;
        RECT 140.460 19.940 145.060 20.110 ;
        RECT 140.460 19.630 140.630 19.940 ;
        RECT 144.890 19.630 145.060 19.940 ;
        RECT 140.430 15.760 140.660 19.630 ;
        RECT 141.260 19.430 144.260 19.600 ;
        RECT 141.030 16.175 141.200 19.215 ;
        RECT 144.320 16.175 144.490 19.215 ;
        RECT 141.260 15.790 144.260 15.960 ;
        RECT 144.870 15.760 145.080 19.630 ;
        RECT 147.010 17.180 147.180 28.670 ;
        RECT 147.490 28.650 149.430 28.670 ;
        RECT 147.810 28.160 149.110 28.330 ;
        RECT 147.580 17.905 147.750 27.945 ;
        RECT 149.170 17.905 149.340 27.945 ;
        RECT 147.810 17.520 149.110 17.690 ;
        RECT 149.740 17.180 149.910 28.670 ;
        RECT 147.010 17.010 149.910 17.180 ;
        RECT 132.130 15.270 138.730 15.440 ;
        RECT 140.460 15.450 140.630 15.760 ;
        RECT 144.890 15.450 145.060 15.760 ;
        RECT 140.460 15.280 145.060 15.450 ;
      LAYER mcon ;
        RECT 116.655 29.960 116.825 30.130 ;
        RECT 117.615 29.980 117.785 30.150 ;
        RECT 117.975 29.980 118.145 30.150 ;
        RECT 118.335 29.980 118.505 30.150 ;
        RECT 118.695 29.980 118.865 30.150 ;
        RECT 119.055 29.980 119.225 30.150 ;
        RECT 119.415 29.980 119.585 30.150 ;
        RECT 119.775 29.980 119.945 30.150 ;
        RECT 120.135 29.980 120.305 30.150 ;
        RECT 116.655 29.600 116.825 29.770 ;
        RECT 116.655 29.240 116.825 29.410 ;
        RECT 116.655 28.880 116.825 29.050 ;
        RECT 112.720 28.665 112.890 28.835 ;
        RECT 113.080 28.665 113.250 28.835 ;
        RECT 113.440 28.665 113.610 28.835 ;
        RECT 113.800 28.665 113.970 28.835 ;
        RECT 114.160 28.665 114.330 28.835 ;
        RECT 113.075 28.160 113.245 28.330 ;
        RECT 113.435 28.160 113.605 28.330 ;
        RECT 113.795 28.160 113.965 28.330 ;
        RECT 112.640 27.520 112.810 27.690 ;
        RECT 112.640 27.160 112.810 27.330 ;
        RECT 112.640 26.800 112.810 26.970 ;
        RECT 112.640 26.440 112.810 26.610 ;
        RECT 112.640 26.080 112.810 26.250 ;
        RECT 112.640 25.720 112.810 25.890 ;
        RECT 112.640 25.360 112.810 25.530 ;
        RECT 112.640 25.000 112.810 25.170 ;
        RECT 112.640 24.640 112.810 24.810 ;
        RECT 112.640 24.280 112.810 24.450 ;
        RECT 112.640 23.920 112.810 24.090 ;
        RECT 112.640 23.560 112.810 23.730 ;
        RECT 112.640 23.200 112.810 23.370 ;
        RECT 112.640 22.840 112.810 23.010 ;
        RECT 112.640 22.480 112.810 22.650 ;
        RECT 112.640 22.120 112.810 22.290 ;
        RECT 112.640 21.760 112.810 21.930 ;
        RECT 112.640 21.400 112.810 21.570 ;
        RECT 112.640 21.040 112.810 21.210 ;
        RECT 112.640 20.680 112.810 20.850 ;
        RECT 112.640 20.320 112.810 20.490 ;
        RECT 112.640 19.960 112.810 20.130 ;
        RECT 112.640 19.600 112.810 19.770 ;
        RECT 112.640 19.240 112.810 19.410 ;
        RECT 112.640 18.880 112.810 19.050 ;
        RECT 112.640 18.520 112.810 18.690 ;
        RECT 112.640 18.160 112.810 18.330 ;
        RECT 114.230 27.520 114.400 27.690 ;
        RECT 114.230 27.160 114.400 27.330 ;
        RECT 114.230 26.800 114.400 26.970 ;
        RECT 114.230 26.440 114.400 26.610 ;
        RECT 114.230 26.080 114.400 26.250 ;
        RECT 114.230 25.720 114.400 25.890 ;
        RECT 114.230 25.360 114.400 25.530 ;
        RECT 114.230 25.000 114.400 25.170 ;
        RECT 114.230 24.640 114.400 24.810 ;
        RECT 114.230 24.280 114.400 24.450 ;
        RECT 114.230 23.920 114.400 24.090 ;
        RECT 114.230 23.560 114.400 23.730 ;
        RECT 114.230 23.200 114.400 23.370 ;
        RECT 114.230 22.840 114.400 23.010 ;
        RECT 114.230 22.480 114.400 22.650 ;
        RECT 114.230 22.120 114.400 22.290 ;
        RECT 114.230 21.760 114.400 21.930 ;
        RECT 114.230 21.400 114.400 21.570 ;
        RECT 114.230 21.040 114.400 21.210 ;
        RECT 114.230 20.680 114.400 20.850 ;
        RECT 114.230 20.320 114.400 20.490 ;
        RECT 114.230 19.960 114.400 20.130 ;
        RECT 114.230 19.600 114.400 19.770 ;
        RECT 114.230 19.240 114.400 19.410 ;
        RECT 114.230 18.880 114.400 19.050 ;
        RECT 114.230 18.520 114.400 18.690 ;
        RECT 114.230 18.160 114.400 18.330 ;
        RECT 113.075 17.520 113.245 17.690 ;
        RECT 113.435 17.520 113.605 17.690 ;
        RECT 113.795 17.520 113.965 17.690 ;
        RECT 116.655 28.520 116.825 28.690 ;
        RECT 116.655 28.160 116.825 28.330 ;
        RECT 116.655 27.800 116.825 27.970 ;
        RECT 116.655 27.440 116.825 27.610 ;
        RECT 116.655 27.080 116.825 27.250 ;
        RECT 116.655 26.720 116.825 26.890 ;
        RECT 117.230 29.420 117.400 29.590 ;
        RECT 117.230 29.060 117.400 29.230 ;
        RECT 117.230 28.700 117.400 28.870 ;
        RECT 117.230 28.340 117.400 28.510 ;
        RECT 117.230 27.980 117.400 28.150 ;
        RECT 117.230 27.620 117.400 27.790 ;
        RECT 117.230 27.260 117.400 27.430 ;
        RECT 117.230 26.900 117.400 27.070 ;
        RECT 120.520 29.420 120.690 29.590 ;
        RECT 120.520 29.060 120.690 29.230 ;
        RECT 120.520 28.700 120.690 28.870 ;
        RECT 120.520 28.340 120.690 28.510 ;
        RECT 120.520 27.980 120.690 28.150 ;
        RECT 120.520 27.620 120.690 27.790 ;
        RECT 120.520 27.260 120.690 27.430 ;
        RECT 120.520 26.900 120.690 27.070 ;
        RECT 116.655 26.360 116.825 26.530 ;
        RECT 117.615 26.340 117.785 26.510 ;
        RECT 117.975 26.340 118.145 26.510 ;
        RECT 118.335 26.340 118.505 26.510 ;
        RECT 118.695 26.340 118.865 26.510 ;
        RECT 119.055 26.340 119.225 26.510 ;
        RECT 119.415 26.340 119.585 26.510 ;
        RECT 119.775 26.340 119.945 26.510 ;
        RECT 120.135 26.340 120.305 26.510 ;
        RECT 124.515 29.960 124.685 30.130 ;
        RECT 124.875 29.960 125.045 30.130 ;
        RECT 125.235 29.960 125.405 30.130 ;
        RECT 125.595 29.960 125.765 30.130 ;
        RECT 125.955 29.960 126.125 30.130 ;
        RECT 126.315 29.960 126.485 30.130 ;
        RECT 126.675 29.960 126.845 30.130 ;
        RECT 127.035 29.960 127.205 30.130 ;
        RECT 127.395 29.960 127.565 30.130 ;
        RECT 127.755 29.960 127.925 30.130 ;
        RECT 128.115 29.960 128.285 30.130 ;
        RECT 128.475 29.960 128.645 30.130 ;
        RECT 128.835 29.960 129.005 30.130 ;
        RECT 124.030 29.445 124.200 29.615 ;
        RECT 124.030 29.085 124.200 29.255 ;
        RECT 124.030 28.725 124.200 28.895 ;
        RECT 124.030 28.365 124.200 28.535 ;
        RECT 124.030 28.005 124.200 28.175 ;
        RECT 124.030 27.645 124.200 27.815 ;
        RECT 124.030 27.285 124.200 27.455 ;
        RECT 124.030 26.925 124.200 27.095 ;
        RECT 129.320 29.445 129.490 29.615 ;
        RECT 129.320 29.085 129.490 29.255 ;
        RECT 129.320 28.725 129.490 28.895 ;
        RECT 129.320 28.365 129.490 28.535 ;
        RECT 129.320 28.005 129.490 28.175 ;
        RECT 129.320 27.645 129.490 27.815 ;
        RECT 129.320 27.285 129.490 27.455 ;
        RECT 129.320 26.925 129.490 27.095 ;
        RECT 124.515 26.410 124.685 26.580 ;
        RECT 124.875 26.410 125.045 26.580 ;
        RECT 125.235 26.410 125.405 26.580 ;
        RECT 125.595 26.410 125.765 26.580 ;
        RECT 125.955 26.410 126.125 26.580 ;
        RECT 126.315 26.410 126.485 26.580 ;
        RECT 126.675 26.410 126.845 26.580 ;
        RECT 127.035 26.410 127.205 26.580 ;
        RECT 127.395 26.410 127.565 26.580 ;
        RECT 127.755 26.410 127.925 26.580 ;
        RECT 128.115 26.410 128.285 26.580 ;
        RECT 128.475 26.410 128.645 26.580 ;
        RECT 128.835 26.410 129.005 26.580 ;
        RECT 132.145 29.820 132.315 29.990 ;
        RECT 133.205 29.840 133.375 30.010 ;
        RECT 133.565 29.840 133.735 30.010 ;
        RECT 133.925 29.840 134.095 30.010 ;
        RECT 134.285 29.840 134.455 30.010 ;
        RECT 134.645 29.840 134.815 30.010 ;
        RECT 135.005 29.840 135.175 30.010 ;
        RECT 135.365 29.840 135.535 30.010 ;
        RECT 135.725 29.840 135.895 30.010 ;
        RECT 136.085 29.840 136.255 30.010 ;
        RECT 136.445 29.840 136.615 30.010 ;
        RECT 136.805 29.840 136.975 30.010 ;
        RECT 137.165 29.840 137.335 30.010 ;
        RECT 137.525 29.840 137.695 30.010 ;
        RECT 138.585 29.820 138.755 29.990 ;
        RECT 132.145 29.460 132.315 29.630 ;
        RECT 132.145 29.100 132.315 29.270 ;
        RECT 132.720 29.280 132.890 29.450 ;
        RECT 138.010 29.280 138.180 29.450 ;
        RECT 138.585 29.460 138.755 29.630 ;
        RECT 138.585 29.100 138.755 29.270 ;
        RECT 132.145 28.740 132.315 28.910 ;
        RECT 133.205 28.720 133.375 28.890 ;
        RECT 133.565 28.720 133.735 28.890 ;
        RECT 133.925 28.720 134.095 28.890 ;
        RECT 134.285 28.720 134.455 28.890 ;
        RECT 134.645 28.720 134.815 28.890 ;
        RECT 135.005 28.720 135.175 28.890 ;
        RECT 135.365 28.720 135.535 28.890 ;
        RECT 135.725 28.720 135.895 28.890 ;
        RECT 136.085 28.720 136.255 28.890 ;
        RECT 136.445 28.720 136.615 28.890 ;
        RECT 136.805 28.720 136.975 28.890 ;
        RECT 137.165 28.720 137.335 28.890 ;
        RECT 137.525 28.720 137.695 28.890 ;
        RECT 138.585 28.740 138.755 28.910 ;
        RECT 141.425 29.980 141.595 30.150 ;
        RECT 141.785 29.980 141.955 30.150 ;
        RECT 142.145 29.980 142.315 30.150 ;
        RECT 142.505 29.980 142.675 30.150 ;
        RECT 142.865 29.980 143.035 30.150 ;
        RECT 143.225 29.980 143.395 30.150 ;
        RECT 143.585 29.980 143.755 30.150 ;
        RECT 143.945 29.980 144.115 30.150 ;
        RECT 144.900 29.900 145.070 30.070 ;
        RECT 141.040 29.360 141.210 29.530 ;
        RECT 144.330 29.360 144.500 29.530 ;
        RECT 144.900 29.540 145.070 29.710 ;
        RECT 144.900 29.180 145.070 29.350 ;
        RECT 141.425 28.740 141.595 28.910 ;
        RECT 141.785 28.740 141.955 28.910 ;
        RECT 142.145 28.740 142.315 28.910 ;
        RECT 142.505 28.740 142.675 28.910 ;
        RECT 142.865 28.740 143.035 28.910 ;
        RECT 143.225 28.740 143.395 28.910 ;
        RECT 143.585 28.740 143.755 28.910 ;
        RECT 143.945 28.740 144.115 28.910 ;
        RECT 144.900 28.820 145.070 28.990 ;
        RECT 147.655 28.670 147.825 28.840 ;
        RECT 148.015 28.670 148.185 28.840 ;
        RECT 148.375 28.670 148.545 28.840 ;
        RECT 148.735 28.670 148.905 28.840 ;
        RECT 149.095 28.670 149.265 28.840 ;
        RECT 140.450 25.880 140.620 26.050 ;
        RECT 141.405 25.900 141.575 26.070 ;
        RECT 141.765 25.900 141.935 26.070 ;
        RECT 142.125 25.900 142.295 26.070 ;
        RECT 142.485 25.900 142.655 26.070 ;
        RECT 142.845 25.900 143.015 26.070 ;
        RECT 143.205 25.900 143.375 26.070 ;
        RECT 143.565 25.900 143.735 26.070 ;
        RECT 143.925 25.900 144.095 26.070 ;
        RECT 140.450 25.520 140.620 25.690 ;
        RECT 144.880 25.880 145.050 26.050 ;
        RECT 140.450 25.160 140.620 25.330 ;
        RECT 140.450 24.800 140.620 24.970 ;
        RECT 140.450 24.440 140.620 24.610 ;
        RECT 140.450 24.080 140.620 24.250 ;
        RECT 140.450 23.720 140.620 23.890 ;
        RECT 116.665 23.495 116.835 23.665 ;
        RECT 117.620 23.515 117.790 23.685 ;
        RECT 117.980 23.515 118.150 23.685 ;
        RECT 118.340 23.515 118.510 23.685 ;
        RECT 118.700 23.515 118.870 23.685 ;
        RECT 119.060 23.515 119.230 23.685 ;
        RECT 119.420 23.515 119.590 23.685 ;
        RECT 119.780 23.515 119.950 23.685 ;
        RECT 120.140 23.515 120.310 23.685 ;
        RECT 116.665 23.135 116.835 23.305 ;
        RECT 121.100 23.495 121.270 23.665 ;
        RECT 116.665 22.775 116.835 22.945 ;
        RECT 116.665 22.415 116.835 22.585 ;
        RECT 116.665 22.055 116.835 22.225 ;
        RECT 116.665 21.695 116.835 21.865 ;
        RECT 116.665 21.335 116.835 21.505 ;
        RECT 116.665 20.975 116.835 21.145 ;
        RECT 116.665 20.615 116.835 20.785 ;
        RECT 116.665 20.255 116.835 20.425 ;
        RECT 117.235 22.955 117.405 23.125 ;
        RECT 117.235 22.595 117.405 22.765 ;
        RECT 117.235 22.235 117.405 22.405 ;
        RECT 117.235 21.875 117.405 22.045 ;
        RECT 117.235 21.515 117.405 21.685 ;
        RECT 117.235 21.155 117.405 21.325 ;
        RECT 117.235 20.795 117.405 20.965 ;
        RECT 117.235 20.435 117.405 20.605 ;
        RECT 120.525 22.955 120.695 23.125 ;
        RECT 120.525 22.595 120.695 22.765 ;
        RECT 120.525 22.235 120.695 22.405 ;
        RECT 120.525 21.875 120.695 22.045 ;
        RECT 120.525 21.515 120.695 21.685 ;
        RECT 120.525 21.155 120.695 21.325 ;
        RECT 120.525 20.795 120.695 20.965 ;
        RECT 120.525 20.435 120.695 20.605 ;
        RECT 121.100 23.135 121.270 23.305 ;
        RECT 121.100 22.775 121.270 22.945 ;
        RECT 121.100 22.415 121.270 22.585 ;
        RECT 140.450 23.360 140.620 23.530 ;
        RECT 140.450 23.000 140.620 23.170 ;
        RECT 140.450 22.640 140.620 22.810 ;
        RECT 141.020 25.340 141.190 25.510 ;
        RECT 141.020 24.980 141.190 25.150 ;
        RECT 141.020 24.620 141.190 24.790 ;
        RECT 141.020 24.260 141.190 24.430 ;
        RECT 141.020 23.900 141.190 24.070 ;
        RECT 141.020 23.540 141.190 23.710 ;
        RECT 141.020 23.180 141.190 23.350 ;
        RECT 141.020 22.820 141.190 22.990 ;
        RECT 144.310 25.340 144.480 25.510 ;
        RECT 144.310 24.980 144.480 25.150 ;
        RECT 144.310 24.620 144.480 24.790 ;
        RECT 144.310 24.260 144.480 24.430 ;
        RECT 144.310 23.900 144.480 24.070 ;
        RECT 144.310 23.540 144.480 23.710 ;
        RECT 144.310 23.180 144.480 23.350 ;
        RECT 144.310 22.820 144.480 22.990 ;
        RECT 144.880 25.520 145.050 25.690 ;
        RECT 144.880 25.160 145.050 25.330 ;
        RECT 144.880 24.800 145.050 24.970 ;
        RECT 144.880 24.440 145.050 24.610 ;
        RECT 144.880 24.080 145.050 24.250 ;
        RECT 144.880 23.720 145.050 23.890 ;
        RECT 144.880 23.360 145.050 23.530 ;
        RECT 144.880 23.000 145.050 23.170 ;
        RECT 140.450 22.280 140.620 22.450 ;
        RECT 144.880 22.640 145.050 22.810 ;
        RECT 141.405 22.260 141.575 22.430 ;
        RECT 141.765 22.260 141.935 22.430 ;
        RECT 142.125 22.260 142.295 22.430 ;
        RECT 142.485 22.260 142.655 22.430 ;
        RECT 142.845 22.260 143.015 22.430 ;
        RECT 143.205 22.260 143.375 22.430 ;
        RECT 143.565 22.260 143.735 22.430 ;
        RECT 143.925 22.260 144.095 22.430 ;
        RECT 144.880 22.280 145.050 22.450 ;
        RECT 121.100 22.055 121.270 22.225 ;
        RECT 121.100 21.695 121.270 21.865 ;
        RECT 121.100 21.335 121.270 21.505 ;
        RECT 121.100 20.975 121.270 21.145 ;
        RECT 121.100 20.615 121.270 20.785 ;
        RECT 116.665 19.895 116.835 20.065 ;
        RECT 121.100 20.255 121.270 20.425 ;
        RECT 117.620 19.875 117.790 20.045 ;
        RECT 117.980 19.875 118.150 20.045 ;
        RECT 118.340 19.875 118.510 20.045 ;
        RECT 118.700 19.875 118.870 20.045 ;
        RECT 119.060 19.875 119.230 20.045 ;
        RECT 119.420 19.875 119.590 20.045 ;
        RECT 119.780 19.875 119.950 20.045 ;
        RECT 120.140 19.875 120.310 20.045 ;
        RECT 121.100 19.895 121.270 20.065 ;
        RECT 132.135 19.355 132.305 19.525 ;
        RECT 133.185 19.330 133.355 19.500 ;
        RECT 133.545 19.330 133.715 19.500 ;
        RECT 133.905 19.330 134.075 19.500 ;
        RECT 134.265 19.330 134.435 19.500 ;
        RECT 134.625 19.330 134.795 19.500 ;
        RECT 134.985 19.330 135.155 19.500 ;
        RECT 135.345 19.330 135.515 19.500 ;
        RECT 135.705 19.330 135.875 19.500 ;
        RECT 136.065 19.330 136.235 19.500 ;
        RECT 136.425 19.330 136.595 19.500 ;
        RECT 136.785 19.330 136.955 19.500 ;
        RECT 137.145 19.330 137.315 19.500 ;
        RECT 137.505 19.330 137.675 19.500 ;
        RECT 132.135 18.995 132.305 19.165 ;
        RECT 132.135 18.635 132.305 18.805 ;
        RECT 132.135 18.275 132.305 18.445 ;
        RECT 132.135 17.915 132.305 18.085 ;
        RECT 116.655 16.960 116.825 17.130 ;
        RECT 117.605 17.040 117.775 17.210 ;
        RECT 117.965 17.040 118.135 17.210 ;
        RECT 118.325 17.040 118.495 17.210 ;
        RECT 118.685 17.040 118.855 17.210 ;
        RECT 119.045 17.040 119.215 17.210 ;
        RECT 119.405 17.040 119.575 17.210 ;
        RECT 119.765 17.040 119.935 17.210 ;
        RECT 120.125 17.040 120.295 17.210 ;
        RECT 121.085 16.960 121.255 17.130 ;
        RECT 132.135 17.555 132.305 17.725 ;
        RECT 132.135 17.195 132.305 17.365 ;
        RECT 116.655 16.600 116.825 16.770 ;
        RECT 116.655 16.240 116.825 16.410 ;
        RECT 117.220 16.420 117.390 16.590 ;
        RECT 120.510 16.420 120.680 16.590 ;
        RECT 121.085 16.600 121.255 16.770 ;
        RECT 121.085 16.240 121.255 16.410 ;
        RECT 116.655 15.880 116.825 16.050 ;
        RECT 117.605 15.800 117.775 15.970 ;
        RECT 117.965 15.800 118.135 15.970 ;
        RECT 118.325 15.800 118.495 15.970 ;
        RECT 118.685 15.800 118.855 15.970 ;
        RECT 119.045 15.800 119.215 15.970 ;
        RECT 119.405 15.800 119.575 15.970 ;
        RECT 119.765 15.800 119.935 15.970 ;
        RECT 120.125 15.800 120.295 15.970 ;
        RECT 121.085 15.880 121.255 16.050 ;
        RECT 123.105 16.890 123.275 17.060 ;
        RECT 124.165 16.910 124.335 17.080 ;
        RECT 124.525 16.910 124.695 17.080 ;
        RECT 124.885 16.910 125.055 17.080 ;
        RECT 125.245 16.910 125.415 17.080 ;
        RECT 125.605 16.910 125.775 17.080 ;
        RECT 125.965 16.910 126.135 17.080 ;
        RECT 126.325 16.910 126.495 17.080 ;
        RECT 126.685 16.910 126.855 17.080 ;
        RECT 127.045 16.910 127.215 17.080 ;
        RECT 127.405 16.910 127.575 17.080 ;
        RECT 127.765 16.910 127.935 17.080 ;
        RECT 128.125 16.910 128.295 17.080 ;
        RECT 128.485 16.910 128.655 17.080 ;
        RECT 129.545 16.890 129.715 17.060 ;
        RECT 123.105 16.530 123.275 16.700 ;
        RECT 123.105 16.170 123.275 16.340 ;
        RECT 123.680 16.350 123.850 16.520 ;
        RECT 128.970 16.350 129.140 16.520 ;
        RECT 129.545 16.530 129.715 16.700 ;
        RECT 129.545 16.170 129.715 16.340 ;
        RECT 123.105 15.810 123.275 15.980 ;
        RECT 124.165 15.790 124.335 15.960 ;
        RECT 124.525 15.790 124.695 15.960 ;
        RECT 124.885 15.790 125.055 15.960 ;
        RECT 125.245 15.790 125.415 15.960 ;
        RECT 125.605 15.790 125.775 15.960 ;
        RECT 125.965 15.790 126.135 15.960 ;
        RECT 126.325 15.790 126.495 15.960 ;
        RECT 126.685 15.790 126.855 15.960 ;
        RECT 127.045 15.790 127.215 15.960 ;
        RECT 127.405 15.790 127.575 15.960 ;
        RECT 127.765 15.790 127.935 15.960 ;
        RECT 128.125 15.790 128.295 15.960 ;
        RECT 128.485 15.790 128.655 15.960 ;
        RECT 129.545 15.810 129.715 15.980 ;
        RECT 132.135 16.835 132.305 17.005 ;
        RECT 132.135 16.475 132.305 16.645 ;
        RECT 132.135 16.115 132.305 16.285 ;
        RECT 132.700 18.815 132.870 18.985 ;
        RECT 132.700 18.455 132.870 18.625 ;
        RECT 132.700 18.095 132.870 18.265 ;
        RECT 132.700 17.735 132.870 17.905 ;
        RECT 132.700 17.375 132.870 17.545 ;
        RECT 132.700 17.015 132.870 17.185 ;
        RECT 132.700 16.655 132.870 16.825 ;
        RECT 132.700 16.295 132.870 16.465 ;
        RECT 137.990 18.815 138.160 18.985 ;
        RECT 137.990 18.455 138.160 18.625 ;
        RECT 137.990 18.095 138.160 18.265 ;
        RECT 137.990 17.735 138.160 17.905 ;
        RECT 137.990 17.375 138.160 17.545 ;
        RECT 137.990 17.015 138.160 17.185 ;
        RECT 137.990 16.655 138.160 16.825 ;
        RECT 137.990 16.295 138.160 16.465 ;
        RECT 132.135 15.755 132.305 15.925 ;
        RECT 133.185 15.780 133.355 15.950 ;
        RECT 133.545 15.780 133.715 15.950 ;
        RECT 133.905 15.780 134.075 15.950 ;
        RECT 134.265 15.780 134.435 15.950 ;
        RECT 134.625 15.780 134.795 15.950 ;
        RECT 134.985 15.780 135.155 15.950 ;
        RECT 135.345 15.780 135.515 15.950 ;
        RECT 135.705 15.780 135.875 15.950 ;
        RECT 136.065 15.780 136.235 15.950 ;
        RECT 136.425 15.780 136.595 15.950 ;
        RECT 136.785 15.780 136.955 15.950 ;
        RECT 137.145 15.780 137.315 15.950 ;
        RECT 137.505 15.780 137.675 15.950 ;
        RECT 140.460 19.410 140.630 19.580 ;
        RECT 141.415 19.430 141.585 19.600 ;
        RECT 141.775 19.430 141.945 19.600 ;
        RECT 142.135 19.430 142.305 19.600 ;
        RECT 142.495 19.430 142.665 19.600 ;
        RECT 142.855 19.430 143.025 19.600 ;
        RECT 143.215 19.430 143.385 19.600 ;
        RECT 143.575 19.430 143.745 19.600 ;
        RECT 143.935 19.430 144.105 19.600 ;
        RECT 140.460 19.050 140.630 19.220 ;
        RECT 144.890 19.410 145.060 19.580 ;
        RECT 140.460 18.690 140.630 18.860 ;
        RECT 140.460 18.330 140.630 18.500 ;
        RECT 140.460 17.970 140.630 18.140 ;
        RECT 140.460 17.610 140.630 17.780 ;
        RECT 140.460 17.250 140.630 17.420 ;
        RECT 140.460 16.890 140.630 17.060 ;
        RECT 140.460 16.530 140.630 16.700 ;
        RECT 140.460 16.170 140.630 16.340 ;
        RECT 141.030 18.870 141.200 19.040 ;
        RECT 141.030 18.510 141.200 18.680 ;
        RECT 141.030 18.150 141.200 18.320 ;
        RECT 141.030 17.790 141.200 17.960 ;
        RECT 141.030 17.430 141.200 17.600 ;
        RECT 141.030 17.070 141.200 17.240 ;
        RECT 141.030 16.710 141.200 16.880 ;
        RECT 141.030 16.350 141.200 16.520 ;
        RECT 144.320 18.870 144.490 19.040 ;
        RECT 144.320 18.510 144.490 18.680 ;
        RECT 144.320 18.150 144.490 18.320 ;
        RECT 144.320 17.790 144.490 17.960 ;
        RECT 144.320 17.430 144.490 17.600 ;
        RECT 144.320 17.070 144.490 17.240 ;
        RECT 144.320 16.710 144.490 16.880 ;
        RECT 144.320 16.350 144.490 16.520 ;
        RECT 144.890 19.050 145.060 19.220 ;
        RECT 144.890 18.690 145.060 18.860 ;
        RECT 144.890 18.330 145.060 18.500 ;
        RECT 144.890 17.970 145.060 18.140 ;
        RECT 144.890 17.610 145.060 17.780 ;
        RECT 144.890 17.250 145.060 17.420 ;
        RECT 144.890 16.890 145.060 17.060 ;
        RECT 148.015 28.160 148.185 28.330 ;
        RECT 148.375 28.160 148.545 28.330 ;
        RECT 148.735 28.160 148.905 28.330 ;
        RECT 147.580 27.520 147.750 27.690 ;
        RECT 147.580 27.160 147.750 27.330 ;
        RECT 147.580 26.800 147.750 26.970 ;
        RECT 147.580 26.440 147.750 26.610 ;
        RECT 147.580 26.080 147.750 26.250 ;
        RECT 147.580 25.720 147.750 25.890 ;
        RECT 147.580 25.360 147.750 25.530 ;
        RECT 147.580 25.000 147.750 25.170 ;
        RECT 147.580 24.640 147.750 24.810 ;
        RECT 147.580 24.280 147.750 24.450 ;
        RECT 147.580 23.920 147.750 24.090 ;
        RECT 147.580 23.560 147.750 23.730 ;
        RECT 147.580 23.200 147.750 23.370 ;
        RECT 147.580 22.840 147.750 23.010 ;
        RECT 147.580 22.480 147.750 22.650 ;
        RECT 147.580 22.120 147.750 22.290 ;
        RECT 147.580 21.760 147.750 21.930 ;
        RECT 147.580 21.400 147.750 21.570 ;
        RECT 147.580 21.040 147.750 21.210 ;
        RECT 147.580 20.680 147.750 20.850 ;
        RECT 147.580 20.320 147.750 20.490 ;
        RECT 147.580 19.960 147.750 20.130 ;
        RECT 147.580 19.600 147.750 19.770 ;
        RECT 147.580 19.240 147.750 19.410 ;
        RECT 147.580 18.880 147.750 19.050 ;
        RECT 147.580 18.520 147.750 18.690 ;
        RECT 147.580 18.160 147.750 18.330 ;
        RECT 149.170 27.520 149.340 27.690 ;
        RECT 149.170 27.160 149.340 27.330 ;
        RECT 149.170 26.800 149.340 26.970 ;
        RECT 149.170 26.440 149.340 26.610 ;
        RECT 149.170 26.080 149.340 26.250 ;
        RECT 149.170 25.720 149.340 25.890 ;
        RECT 149.170 25.360 149.340 25.530 ;
        RECT 149.170 25.000 149.340 25.170 ;
        RECT 149.170 24.640 149.340 24.810 ;
        RECT 149.170 24.280 149.340 24.450 ;
        RECT 149.170 23.920 149.340 24.090 ;
        RECT 149.170 23.560 149.340 23.730 ;
        RECT 149.170 23.200 149.340 23.370 ;
        RECT 149.170 22.840 149.340 23.010 ;
        RECT 149.170 22.480 149.340 22.650 ;
        RECT 149.170 22.120 149.340 22.290 ;
        RECT 149.170 21.760 149.340 21.930 ;
        RECT 149.170 21.400 149.340 21.570 ;
        RECT 149.170 21.040 149.340 21.210 ;
        RECT 149.170 20.680 149.340 20.850 ;
        RECT 149.170 20.320 149.340 20.490 ;
        RECT 149.170 19.960 149.340 20.130 ;
        RECT 149.170 19.600 149.340 19.770 ;
        RECT 149.170 19.240 149.340 19.410 ;
        RECT 149.170 18.880 149.340 19.050 ;
        RECT 149.170 18.520 149.340 18.690 ;
        RECT 149.170 18.160 149.340 18.330 ;
        RECT 148.015 17.520 148.185 17.690 ;
        RECT 148.375 17.520 148.545 17.690 ;
        RECT 148.735 17.520 148.905 17.690 ;
        RECT 144.890 16.530 145.060 16.700 ;
        RECT 140.460 15.810 140.630 15.980 ;
        RECT 144.890 16.170 145.060 16.340 ;
        RECT 141.415 15.790 141.585 15.960 ;
        RECT 141.775 15.790 141.945 15.960 ;
        RECT 142.135 15.790 142.305 15.960 ;
        RECT 142.495 15.790 142.665 15.960 ;
        RECT 142.855 15.790 143.025 15.960 ;
        RECT 143.215 15.790 143.385 15.960 ;
        RECT 143.575 15.790 143.745 15.960 ;
        RECT 143.935 15.790 144.105 15.960 ;
        RECT 144.890 15.810 145.060 15.980 ;
      LAYER met1 ;
        RECT 151.020 34.210 152.020 34.240 ;
        RECT 106.040 32.530 109.030 33.350 ;
        RECT 113.090 33.210 152.020 34.210 ;
        RECT 151.020 33.180 152.020 33.210 ;
        RECT 106.040 32.000 150.080 32.530 ;
        RECT 106.040 31.730 109.030 32.000 ;
        RECT 113.120 28.960 114.120 31.710 ;
        RECT 116.630 30.720 116.870 32.000 ;
        RECT 138.080 31.180 141.140 31.370 ;
        RECT 111.970 28.580 115.080 28.960 ;
        RECT 116.570 28.370 116.920 30.720 ;
        RECT 117.480 29.950 120.440 30.180 ;
        RECT 124.280 29.930 129.240 30.160 ;
        RECT 117.200 28.370 117.430 29.745 ;
        RECT 112.890 28.340 114.150 28.360 ;
        RECT 112.630 28.130 114.150 28.340 ;
        RECT 116.570 28.140 117.430 28.370 ;
        RECT 112.630 27.925 112.930 28.130 ;
        RECT 112.610 27.900 112.930 27.925 ;
        RECT 112.610 18.080 112.840 27.900 ;
        RECT 112.540 17.925 112.840 18.080 ;
        RECT 114.200 18.550 114.430 27.925 ;
        RECT 116.570 21.870 116.920 28.140 ;
        RECT 117.200 26.745 117.430 28.140 ;
        RECT 120.490 28.430 120.720 29.745 ;
        RECT 120.490 28.170 123.330 28.430 ;
        RECT 120.490 26.745 120.720 28.170 ;
        RECT 124.000 26.770 124.230 29.770 ;
        RECT 129.290 26.770 129.520 29.770 ;
        RECT 132.060 29.460 132.410 30.600 ;
        RECT 132.970 29.810 137.930 30.040 ;
        RECT 138.080 29.650 138.300 31.180 ;
        RECT 132.690 29.460 132.920 29.650 ;
        RECT 130.190 29.150 132.920 29.460 ;
        RECT 132.060 28.140 132.410 29.150 ;
        RECT 132.690 29.080 132.920 29.150 ;
        RECT 137.980 29.560 138.300 29.650 ;
        RECT 137.980 29.080 138.210 29.560 ;
        RECT 133.150 28.920 133.510 28.950 ;
        RECT 132.970 28.690 137.930 28.920 ;
        RECT 117.480 26.310 120.440 26.540 ;
        RECT 124.280 26.380 129.240 26.610 ;
        RECT 118.750 23.715 119.050 26.310 ;
        RECT 128.710 25.190 129.050 25.770 ;
        RECT 133.150 25.190 133.510 28.690 ;
        RECT 138.490 28.130 138.870 30.610 ;
        RECT 140.920 29.745 141.140 31.180 ;
        RECT 144.900 30.740 145.140 32.000 ;
        RECT 150.700 30.810 151.700 30.840 ;
        RECT 141.290 29.950 144.250 30.180 ;
        RECT 140.920 29.560 141.240 29.745 ;
        RECT 141.010 29.460 141.240 29.560 ;
        RECT 144.300 29.510 144.530 29.745 ;
        RECT 144.810 29.510 145.180 30.740 ;
        RECT 148.365 29.810 151.700 30.810 ;
        RECT 141.010 29.200 141.250 29.460 ;
        RECT 144.300 29.300 145.180 29.510 ;
        RECT 141.010 29.145 141.240 29.200 ;
        RECT 144.300 29.145 144.530 29.300 ;
        RECT 141.290 28.710 144.250 28.940 ;
        RECT 128.710 24.820 133.510 25.190 ;
        RECT 128.710 24.810 129.050 24.820 ;
        RECT 117.485 23.700 120.445 23.715 ;
        RECT 117.485 23.485 120.710 23.700 ;
        RECT 120.380 23.280 120.710 23.485 ;
        RECT 117.205 21.870 117.435 23.280 ;
        RECT 120.380 23.040 120.725 23.280 ;
        RECT 116.570 21.650 117.435 21.870 ;
        RECT 116.570 19.310 116.920 21.650 ;
        RECT 117.205 20.280 117.435 21.650 ;
        RECT 120.495 20.280 120.725 23.040 ;
        RECT 117.485 19.845 120.445 20.075 ;
        RECT 118.750 18.550 119.050 19.845 ;
        RECT 114.200 18.290 119.050 18.550 ;
        RECT 114.200 17.925 114.430 18.290 ;
        RECT 104.000 14.030 109.020 14.830 ;
        RECT 112.540 14.030 112.740 17.925 ;
        RECT 112.890 17.490 114.150 17.720 ;
        RECT 116.570 16.610 116.920 17.770 ;
        RECT 118.750 17.240 119.050 18.290 ;
        RECT 117.470 17.010 120.430 17.240 ;
        RECT 117.190 16.610 117.420 16.805 ;
        RECT 116.570 16.400 117.420 16.610 ;
        RECT 116.570 15.250 116.920 16.400 ;
        RECT 117.190 16.205 117.420 16.400 ;
        RECT 120.480 16.510 120.710 16.805 ;
        RECT 120.480 16.205 120.820 16.510 ;
        RECT 117.470 15.770 120.430 16.000 ;
        RECT 120.580 14.940 120.820 16.205 ;
        RECT 121.020 15.200 121.340 24.310 ;
        RECT 138.540 23.120 138.810 28.130 ;
        RECT 123.030 22.780 138.810 23.120 ;
        RECT 123.030 17.670 123.350 22.780 ;
        RECT 128.650 20.740 133.450 21.110 ;
        RECT 122.980 15.210 123.370 17.670 ;
        RECT 128.650 17.110 129.010 20.740 ;
        RECT 123.930 16.980 129.010 17.110 ;
        RECT 123.930 16.880 128.890 16.980 ;
        RECT 123.650 16.510 123.880 16.720 ;
        RECT 123.530 16.150 123.880 16.510 ;
        RECT 128.940 16.620 129.170 16.720 ;
        RECT 129.470 16.620 129.840 17.670 ;
        RECT 132.050 16.620 132.370 20.120 ;
        RECT 133.110 19.530 133.450 20.740 ;
        RECT 132.950 19.520 137.910 19.530 ;
        RECT 132.950 19.300 138.150 19.520 ;
        RECT 137.810 19.140 138.150 19.300 ;
        RECT 132.670 16.620 132.900 19.140 ;
        RECT 137.810 19.030 138.190 19.140 ;
        RECT 128.940 16.310 132.900 16.620 ;
        RECT 128.940 16.150 129.170 16.310 ;
        RECT 121.700 14.940 122.660 15.210 ;
        RECT 123.530 14.940 123.770 16.150 ;
        RECT 123.930 15.760 128.890 15.990 ;
        RECT 129.470 15.200 129.840 16.310 ;
        RECT 120.580 14.680 123.770 14.940 ;
        RECT 121.700 14.250 122.660 14.680 ;
        RECT 130.570 14.030 131.030 16.310 ;
        RECT 132.050 15.210 132.370 16.310 ;
        RECT 132.670 16.140 132.900 16.310 ;
        RECT 137.960 16.390 138.190 19.030 ;
        RECT 137.960 16.140 138.370 16.390 ;
        RECT 132.950 15.750 137.910 15.980 ;
        RECT 138.150 14.920 138.370 16.140 ;
        RECT 140.370 15.200 140.730 26.680 ;
        RECT 142.460 26.100 142.760 28.710 ;
        RECT 141.270 25.870 144.230 26.100 ;
        RECT 140.990 22.940 141.220 25.665 ;
        RECT 144.280 24.240 144.510 25.665 ;
        RECT 144.810 24.240 145.180 29.300 ;
        RECT 148.385 28.930 149.350 29.810 ;
        RECT 150.700 29.780 151.700 29.810 ;
        RECT 146.950 28.590 150.000 28.930 ;
        RECT 147.830 28.310 149.090 28.360 ;
        RECT 147.830 28.130 149.360 28.310 ;
        RECT 149.060 27.925 149.360 28.130 ;
        RECT 144.280 24.040 145.180 24.240 ;
        RECT 140.990 22.665 141.360 22.940 ;
        RECT 144.280 22.665 144.510 24.040 ;
        RECT 141.030 22.460 141.360 22.665 ;
        RECT 141.030 22.280 144.230 22.460 ;
        RECT 141.270 22.230 144.230 22.280 ;
        RECT 142.810 20.960 143.110 22.230 ;
        RECT 144.810 21.660 145.180 24.040 ;
        RECT 147.550 20.960 147.780 27.925 ;
        RECT 149.060 27.870 149.370 27.925 ;
        RECT 142.810 20.700 147.780 20.960 ;
        RECT 142.810 19.630 143.110 20.700 ;
        RECT 141.280 19.400 144.240 19.630 ;
        RECT 141.000 16.390 141.230 19.195 ;
        RECT 140.910 16.195 141.230 16.390 ;
        RECT 144.290 17.790 144.520 19.195 ;
        RECT 144.820 17.790 145.160 20.190 ;
        RECT 147.550 17.925 147.780 20.700 ;
        RECT 149.140 18.090 149.370 27.870 ;
        RECT 149.140 17.925 149.460 18.090 ;
        RECT 144.290 17.590 145.160 17.790 ;
        RECT 144.290 16.195 144.520 17.590 ;
        RECT 140.910 14.920 141.130 16.195 ;
        RECT 141.280 15.760 144.240 15.990 ;
        RECT 144.820 15.190 145.160 17.590 ;
        RECT 147.830 17.490 149.090 17.720 ;
        RECT 138.150 14.660 141.130 14.920 ;
        RECT 149.260 14.030 149.460 17.925 ;
        RECT 104.000 13.500 150.080 14.030 ;
        RECT 104.000 13.210 109.020 13.500 ;
      LAYER via ;
        RECT 106.080 31.730 107.700 33.350 ;
        RECT 113.120 33.210 114.120 34.210 ;
        RECT 151.020 33.210 152.020 34.210 ;
        RECT 113.120 30.680 114.120 31.680 ;
        RECT 150.700 29.810 151.700 30.810 ;
        RECT 104.040 13.210 105.660 14.830 ;
        RECT 121.730 14.280 122.630 15.180 ;
      LAYER met2 ;
        RECT 102.990 31.730 107.730 33.350 ;
        RECT 113.120 30.650 114.120 34.240 ;
        RECT 150.990 34.190 152.050 34.210 ;
        RECT 150.990 33.230 153.790 34.190 ;
        RECT 150.990 33.210 152.050 33.230 ;
        RECT 150.670 30.790 151.730 30.810 ;
        RECT 150.670 29.830 153.470 30.790 ;
        RECT 150.670 29.810 151.730 29.830 ;
        RECT 100.950 13.210 105.690 14.830 ;
        RECT 121.730 12.280 122.630 15.210 ;
      LAYER via2 ;
        RECT 103.040 31.770 104.580 33.310 ;
        RECT 152.780 33.230 153.740 34.190 ;
        RECT 152.460 29.830 153.420 30.790 ;
        RECT 101.000 13.250 102.540 14.790 ;
        RECT 121.755 12.325 122.605 13.175 ;
      LAYER met3 ;
        RECT 152.755 34.170 153.765 34.215 ;
        RECT 37.285 33.320 38.835 33.345 ;
        RECT 37.280 31.760 61.280 33.320 ;
        RECT 103.015 33.310 104.605 33.335 ;
        RECT 99.400 31.770 104.605 33.310 ;
        RECT 152.755 33.250 155.690 34.170 ;
        RECT 152.755 33.205 153.765 33.250 ;
        RECT 37.285 31.735 38.835 31.760 ;
        RECT 103.015 31.745 104.605 31.770 ;
        RECT 152.435 30.770 153.445 30.815 ;
        RECT 152.435 29.850 155.370 30.770 ;
        RECT 152.435 29.805 153.445 29.850 ;
        RECT 100.975 14.790 102.565 14.815 ;
        RECT 97.360 13.250 102.565 14.790 ;
        RECT 100.975 13.225 102.565 13.250 ;
        RECT 121.730 11.720 122.630 13.200 ;
        RECT 121.700 10.820 122.660 11.720 ;
      LAYER via3 ;
        RECT 37.285 31.765 38.835 33.315 ;
        RECT 59.695 31.765 61.245 33.315 ;
        RECT 99.435 31.775 100.965 33.305 ;
        RECT 154.740 33.250 155.660 34.170 ;
        RECT 154.420 29.850 155.340 30.770 ;
        RECT 97.395 13.255 98.925 14.785 ;
        RECT 121.730 10.820 122.630 11.720 ;
      LAYER met4 ;
        RECT 3.990 223.710 4.290 224.760 ;
        RECT 7.670 223.710 7.970 224.760 ;
        RECT 11.350 223.710 11.650 224.760 ;
        RECT 15.030 223.710 15.330 224.760 ;
        RECT 18.710 223.710 19.010 224.760 ;
        RECT 22.390 223.710 22.690 224.760 ;
        RECT 26.070 223.710 26.370 224.760 ;
        RECT 29.750 223.710 30.050 224.760 ;
        RECT 33.430 223.710 33.730 224.760 ;
        RECT 37.110 223.710 37.410 224.760 ;
        RECT 40.790 223.710 41.090 224.760 ;
        RECT 44.470 223.710 44.770 224.760 ;
        RECT 48.150 223.710 48.450 224.760 ;
        RECT 51.830 223.710 52.130 224.760 ;
        RECT 55.510 223.710 55.810 224.760 ;
        RECT 59.190 223.710 59.490 224.760 ;
        RECT 62.870 223.710 63.170 224.760 ;
        RECT 66.550 223.710 66.850 224.760 ;
        RECT 70.230 223.710 70.530 224.760 ;
        RECT 73.910 223.710 74.210 224.760 ;
        RECT 77.590 223.710 77.890 224.760 ;
        RECT 81.270 223.710 81.570 224.760 ;
        RECT 84.950 223.710 85.250 224.760 ;
        RECT 88.630 223.710 88.930 224.760 ;
        RECT 3.990 223.410 88.930 223.710 ;
        RECT 49.000 220.760 50.500 223.410 ;
        RECT 154.735 34.160 155.665 34.175 ;
        RECT 37.280 33.290 38.840 33.320 ;
        RECT 2.500 31.790 38.840 33.290 ;
        RECT 37.280 31.760 38.840 31.790 ;
        RECT 59.690 33.290 61.250 33.320 ;
        RECT 99.430 33.290 100.970 33.310 ;
        RECT 59.690 31.790 100.970 33.290 ;
        RECT 154.735 33.260 157.310 34.160 ;
        RECT 154.735 33.245 155.665 33.260 ;
        RECT 59.690 31.760 61.250 31.790 ;
        RECT 99.430 31.770 100.970 31.790 ;
        RECT 154.415 30.760 155.345 30.775 ;
        RECT 154.415 29.860 155.370 30.760 ;
        RECT 154.415 29.845 155.345 29.860 ;
        RECT 97.390 14.770 98.930 14.790 ;
        RECT 50.500 13.270 98.930 14.770 ;
        RECT 97.390 13.250 98.930 13.270 ;
        RECT 121.725 10.815 122.635 11.725 ;
        RECT 121.730 9.580 122.630 10.815 ;
        RECT 112.250 8.680 122.630 9.580 ;
        RECT 154.430 9.530 155.330 29.845 ;
        RECT 112.250 1.000 113.150 8.680 ;
        RECT 134.330 8.630 155.330 9.530 ;
        RECT 134.330 1.000 135.230 8.630 ;
        RECT 156.410 1.000 157.310 33.260 ;
  END
END tt_um_adennen_inverter
END LIBRARY

